  --Example instantiation for system 'nios2'
  nios2_inst : nios2
    port map(
      altpll_0_c0 => altpll_0_c0,
      altpll_0_c1_out => altpll_0_c1_out,
      locked_from_the_altpll_0 => locked_from_the_altpll_0,
      out_port_from_the_cal_dac_code_pio => out_port_from_the_cal_dac_code_pio,
      out_port_from_the_gen_code_strobe => out_port_from_the_gen_code_strobe,
      out_port_from_the_gen_code_value_pio_0 => out_port_from_the_gen_code_value_pio_0,
      out_port_from_the_gen_code_value_pio_1 => out_port_from_the_gen_code_value_pio_1,
      out_port_from_the_latch_pio => out_port_from_the_latch_pio,
      out_port_from_the_led_pio => out_port_from_the_led_pio,
      out_port_from_the_sample_and_hold_pio => out_port_from_the_sample_and_hold_pio,
      out_port_from_the_switch_pio => out_port_from_the_switch_pio,
      out_port_from_the_usb_code_pio => out_port_from_the_usb_code_pio,
      phasedone_from_the_altpll_0 => phasedone_from_the_altpll_0,
      zs_addr_from_the_sdram_0 => zs_addr_from_the_sdram_0,
      zs_ba_from_the_sdram_0 => zs_ba_from_the_sdram_0,
      zs_cas_n_from_the_sdram_0 => zs_cas_n_from_the_sdram_0,
      zs_cke_from_the_sdram_0 => zs_cke_from_the_sdram_0,
      zs_cs_n_from_the_sdram_0 => zs_cs_n_from_the_sdram_0,
      zs_dq_to_and_from_the_sdram_0 => zs_dq_to_and_from_the_sdram_0,
      zs_dqm_from_the_sdram_0 => zs_dqm_from_the_sdram_0,
      zs_ras_n_from_the_sdram_0 => zs_ras_n_from_the_sdram_0,
      zs_we_n_from_the_sdram_0 => zs_we_n_from_the_sdram_0,
      clk_0 => clk_0,
      in_port_to_the_comparator_pio => in_port_to_the_comparator_pio,
      in_port_to_the_mode_select => in_port_to_the_mode_select,
      processor_clk => processor_clk,
      reset_n => reset_n
    );


