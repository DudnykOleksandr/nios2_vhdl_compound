--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2012 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity altpll_0_pll_slave_arbitrator is 
        port (
              -- inputs:
                 signal altpll_0_pll_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_5_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_5_out_read : IN STD_LOGIC;
                 signal nios2_clock_5_out_write : IN STD_LOGIC;
                 signal nios2_clock_5_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal altpll_0_pll_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal altpll_0_pll_slave_read : OUT STD_LOGIC;
                 signal altpll_0_pll_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal altpll_0_pll_slave_reset : OUT STD_LOGIC;
                 signal altpll_0_pll_slave_write : OUT STD_LOGIC;
                 signal altpll_0_pll_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_altpll_0_pll_slave_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_5_out_granted_altpll_0_pll_slave : OUT STD_LOGIC;
                 signal nios2_clock_5_out_qualified_request_altpll_0_pll_slave : OUT STD_LOGIC;
                 signal nios2_clock_5_out_read_data_valid_altpll_0_pll_slave : OUT STD_LOGIC;
                 signal nios2_clock_5_out_requests_altpll_0_pll_slave : OUT STD_LOGIC
              );
end entity altpll_0_pll_slave_arbitrator;


architecture europa of altpll_0_pll_slave_arbitrator is
                signal altpll_0_pll_slave_allgrants :  STD_LOGIC;
                signal altpll_0_pll_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal altpll_0_pll_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal altpll_0_pll_slave_any_continuerequest :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_counter_enable :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_share_counter :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_share_set_values :  STD_LOGIC;
                signal altpll_0_pll_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal altpll_0_pll_slave_begins_xfer :  STD_LOGIC;
                signal altpll_0_pll_slave_end_xfer :  STD_LOGIC;
                signal altpll_0_pll_slave_firsttransfer :  STD_LOGIC;
                signal altpll_0_pll_slave_grant_vector :  STD_LOGIC;
                signal altpll_0_pll_slave_in_a_read_cycle :  STD_LOGIC;
                signal altpll_0_pll_slave_in_a_write_cycle :  STD_LOGIC;
                signal altpll_0_pll_slave_master_qreq_vector :  STD_LOGIC;
                signal altpll_0_pll_slave_non_bursting_master_requests :  STD_LOGIC;
                signal altpll_0_pll_slave_reg_firsttransfer :  STD_LOGIC;
                signal altpll_0_pll_slave_slavearbiterlockenable :  STD_LOGIC;
                signal altpll_0_pll_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal altpll_0_pll_slave_unreg_firsttransfer :  STD_LOGIC;
                signal altpll_0_pll_slave_waits_for_read :  STD_LOGIC;
                signal altpll_0_pll_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_altpll_0_pll_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_5_out_granted_altpll_0_pll_slave :  STD_LOGIC;
                signal internal_nios2_clock_5_out_qualified_request_altpll_0_pll_slave :  STD_LOGIC;
                signal internal_nios2_clock_5_out_requests_altpll_0_pll_slave :  STD_LOGIC;
                signal nios2_clock_5_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_5_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_5_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_5_out_saved_grant_altpll_0_pll_slave :  STD_LOGIC;
                signal shifted_address_to_altpll_0_pll_slave_from_nios2_clock_5_out :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal wait_for_altpll_0_pll_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT altpll_0_pll_slave_end_xfer;
    end if;

  end process;

  altpll_0_pll_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_5_out_qualified_request_altpll_0_pll_slave);
  --assign altpll_0_pll_slave_readdata_from_sa = altpll_0_pll_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  altpll_0_pll_slave_readdata_from_sa <= altpll_0_pll_slave_readdata;
  internal_nios2_clock_5_out_requests_altpll_0_pll_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_5_out_read OR nios2_clock_5_out_write)))))));
  --altpll_0_pll_slave_arb_share_counter set values, which is an e_mux
  altpll_0_pll_slave_arb_share_set_values <= std_logic'('1');
  --altpll_0_pll_slave_non_bursting_master_requests mux, which is an e_mux
  altpll_0_pll_slave_non_bursting_master_requests <= internal_nios2_clock_5_out_requests_altpll_0_pll_slave;
  --altpll_0_pll_slave_any_bursting_master_saved_grant mux, which is an e_mux
  altpll_0_pll_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --altpll_0_pll_slave_arb_share_counter_next_value assignment, which is an e_assign
  altpll_0_pll_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(altpll_0_pll_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(altpll_0_pll_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --altpll_0_pll_slave_allgrants all slave grants, which is an e_mux
  altpll_0_pll_slave_allgrants <= altpll_0_pll_slave_grant_vector;
  --altpll_0_pll_slave_end_xfer assignment, which is an e_assign
  altpll_0_pll_slave_end_xfer <= NOT ((altpll_0_pll_slave_waits_for_read OR altpll_0_pll_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_altpll_0_pll_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_altpll_0_pll_slave <= altpll_0_pll_slave_end_xfer AND (((NOT altpll_0_pll_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --altpll_0_pll_slave_arb_share_counter arbitration counter enable, which is an e_assign
  altpll_0_pll_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_altpll_0_pll_slave AND altpll_0_pll_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_altpll_0_pll_slave AND NOT altpll_0_pll_slave_non_bursting_master_requests));
  --altpll_0_pll_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_0_pll_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(altpll_0_pll_slave_arb_counter_enable) = '1' then 
        altpll_0_pll_slave_arb_share_counter <= altpll_0_pll_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --altpll_0_pll_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_0_pll_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((altpll_0_pll_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_altpll_0_pll_slave)) OR ((end_xfer_arb_share_counter_term_altpll_0_pll_slave AND NOT altpll_0_pll_slave_non_bursting_master_requests)))) = '1' then 
        altpll_0_pll_slave_slavearbiterlockenable <= altpll_0_pll_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_5/out altpll_0/pll_slave arbiterlock, which is an e_assign
  nios2_clock_5_out_arbiterlock <= altpll_0_pll_slave_slavearbiterlockenable AND nios2_clock_5_out_continuerequest;
  --altpll_0_pll_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  altpll_0_pll_slave_slavearbiterlockenable2 <= altpll_0_pll_slave_arb_share_counter_next_value;
  --nios2_clock_5/out altpll_0/pll_slave arbiterlock2, which is an e_assign
  nios2_clock_5_out_arbiterlock2 <= altpll_0_pll_slave_slavearbiterlockenable2 AND nios2_clock_5_out_continuerequest;
  --altpll_0_pll_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  altpll_0_pll_slave_any_continuerequest <= std_logic'('1');
  --nios2_clock_5_out_continuerequest continued request, which is an e_assign
  nios2_clock_5_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_5_out_qualified_request_altpll_0_pll_slave <= internal_nios2_clock_5_out_requests_altpll_0_pll_slave;
  --altpll_0_pll_slave_writedata mux, which is an e_mux
  altpll_0_pll_slave_writedata <= nios2_clock_5_out_writedata;
  --master is always granted when requested
  internal_nios2_clock_5_out_granted_altpll_0_pll_slave <= internal_nios2_clock_5_out_qualified_request_altpll_0_pll_slave;
  --nios2_clock_5/out saved-grant altpll_0/pll_slave, which is an e_assign
  nios2_clock_5_out_saved_grant_altpll_0_pll_slave <= internal_nios2_clock_5_out_requests_altpll_0_pll_slave;
  --allow new arb cycle for altpll_0/pll_slave, which is an e_assign
  altpll_0_pll_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  altpll_0_pll_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  altpll_0_pll_slave_master_qreq_vector <= std_logic'('1');
  --~altpll_0_pll_slave_reset assignment, which is an e_assign
  altpll_0_pll_slave_reset <= NOT reset_n;
  --altpll_0_pll_slave_firsttransfer first transaction, which is an e_assign
  altpll_0_pll_slave_firsttransfer <= A_WE_StdLogic((std_logic'(altpll_0_pll_slave_begins_xfer) = '1'), altpll_0_pll_slave_unreg_firsttransfer, altpll_0_pll_slave_reg_firsttransfer);
  --altpll_0_pll_slave_unreg_firsttransfer first transaction, which is an e_assign
  altpll_0_pll_slave_unreg_firsttransfer <= NOT ((altpll_0_pll_slave_slavearbiterlockenable AND altpll_0_pll_slave_any_continuerequest));
  --altpll_0_pll_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_0_pll_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(altpll_0_pll_slave_begins_xfer) = '1' then 
        altpll_0_pll_slave_reg_firsttransfer <= altpll_0_pll_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --altpll_0_pll_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  altpll_0_pll_slave_beginbursttransfer_internal <= altpll_0_pll_slave_begins_xfer;
  --altpll_0_pll_slave_read assignment, which is an e_mux
  altpll_0_pll_slave_read <= internal_nios2_clock_5_out_granted_altpll_0_pll_slave AND nios2_clock_5_out_read;
  --altpll_0_pll_slave_write assignment, which is an e_mux
  altpll_0_pll_slave_write <= internal_nios2_clock_5_out_granted_altpll_0_pll_slave AND nios2_clock_5_out_write;
  shifted_address_to_altpll_0_pll_slave_from_nios2_clock_5_out <= nios2_clock_5_out_address_to_slave;
  --altpll_0_pll_slave_address mux, which is an e_mux
  altpll_0_pll_slave_address <= A_EXT (A_SRL(shifted_address_to_altpll_0_pll_slave_from_nios2_clock_5_out,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_altpll_0_pll_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_altpll_0_pll_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_altpll_0_pll_slave_end_xfer <= altpll_0_pll_slave_end_xfer;
    end if;

  end process;

  --altpll_0_pll_slave_waits_for_read in a cycle, which is an e_mux
  altpll_0_pll_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --altpll_0_pll_slave_in_a_read_cycle assignment, which is an e_assign
  altpll_0_pll_slave_in_a_read_cycle <= internal_nios2_clock_5_out_granted_altpll_0_pll_slave AND nios2_clock_5_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= altpll_0_pll_slave_in_a_read_cycle;
  --altpll_0_pll_slave_waits_for_write in a cycle, which is an e_mux
  altpll_0_pll_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --altpll_0_pll_slave_in_a_write_cycle assignment, which is an e_assign
  altpll_0_pll_slave_in_a_write_cycle <= internal_nios2_clock_5_out_granted_altpll_0_pll_slave AND nios2_clock_5_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= altpll_0_pll_slave_in_a_write_cycle;
  wait_for_altpll_0_pll_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_5_out_granted_altpll_0_pll_slave <= internal_nios2_clock_5_out_granted_altpll_0_pll_slave;
  --vhdl renameroo for output signals
  nios2_clock_5_out_qualified_request_altpll_0_pll_slave <= internal_nios2_clock_5_out_qualified_request_altpll_0_pll_slave;
  --vhdl renameroo for output signals
  nios2_clock_5_out_requests_altpll_0_pll_slave <= internal_nios2_clock_5_out_requests_altpll_0_pll_slave;
--synthesis translate_off
    --altpll_0/pll_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cal_dac_code_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal cal_dac_code_pio_s1_readdata : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_15_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_15_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_15_out_read : IN STD_LOGIC;
                 signal nios2_clock_15_out_write : IN STD_LOGIC;
                 signal nios2_clock_15_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cal_dac_code_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cal_dac_code_pio_s1_chipselect : OUT STD_LOGIC;
                 signal cal_dac_code_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal cal_dac_code_pio_s1_reset_n : OUT STD_LOGIC;
                 signal cal_dac_code_pio_s1_write_n : OUT STD_LOGIC;
                 signal cal_dac_code_pio_s1_writedata : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal d1_cal_dac_code_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_15_out_granted_cal_dac_code_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_15_out_requests_cal_dac_code_pio_s1 : OUT STD_LOGIC
              );
end entity cal_dac_code_pio_s1_arbitrator;


architecture europa of cal_dac_code_pio_s1_arbitrator is
                signal cal_dac_code_pio_s1_allgrants :  STD_LOGIC;
                signal cal_dac_code_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal cal_dac_code_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cal_dac_code_pio_s1_any_continuerequest :  STD_LOGIC;
                signal cal_dac_code_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal cal_dac_code_pio_s1_arb_share_counter :  STD_LOGIC;
                signal cal_dac_code_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal cal_dac_code_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal cal_dac_code_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal cal_dac_code_pio_s1_begins_xfer :  STD_LOGIC;
                signal cal_dac_code_pio_s1_end_xfer :  STD_LOGIC;
                signal cal_dac_code_pio_s1_firsttransfer :  STD_LOGIC;
                signal cal_dac_code_pio_s1_grant_vector :  STD_LOGIC;
                signal cal_dac_code_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal cal_dac_code_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal cal_dac_code_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal cal_dac_code_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal cal_dac_code_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal cal_dac_code_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal cal_dac_code_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal cal_dac_code_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal cal_dac_code_pio_s1_waits_for_read :  STD_LOGIC;
                signal cal_dac_code_pio_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_15_out_granted_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_15_out_requests_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_15_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_15_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_15_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_15_out_saved_grant_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal wait_for_cal_dac_code_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cal_dac_code_pio_s1_end_xfer;
    end if;

  end process;

  cal_dac_code_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1);
  --assign cal_dac_code_pio_s1_readdata_from_sa = cal_dac_code_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cal_dac_code_pio_s1_readdata_from_sa <= cal_dac_code_pio_s1_readdata;
  internal_nios2_clock_15_out_requests_cal_dac_code_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_15_out_read OR nios2_clock_15_out_write)))))));
  --cal_dac_code_pio_s1_arb_share_counter set values, which is an e_mux
  cal_dac_code_pio_s1_arb_share_set_values <= std_logic'('1');
  --cal_dac_code_pio_s1_non_bursting_master_requests mux, which is an e_mux
  cal_dac_code_pio_s1_non_bursting_master_requests <= internal_nios2_clock_15_out_requests_cal_dac_code_pio_s1;
  --cal_dac_code_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  cal_dac_code_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --cal_dac_code_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  cal_dac_code_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cal_dac_code_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cal_dac_code_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(cal_dac_code_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cal_dac_code_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --cal_dac_code_pio_s1_allgrants all slave grants, which is an e_mux
  cal_dac_code_pio_s1_allgrants <= cal_dac_code_pio_s1_grant_vector;
  --cal_dac_code_pio_s1_end_xfer assignment, which is an e_assign
  cal_dac_code_pio_s1_end_xfer <= NOT ((cal_dac_code_pio_s1_waits_for_read OR cal_dac_code_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_cal_dac_code_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cal_dac_code_pio_s1 <= cal_dac_code_pio_s1_end_xfer AND (((NOT cal_dac_code_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cal_dac_code_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  cal_dac_code_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cal_dac_code_pio_s1 AND cal_dac_code_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_cal_dac_code_pio_s1 AND NOT cal_dac_code_pio_s1_non_bursting_master_requests));
  --cal_dac_code_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cal_dac_code_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(cal_dac_code_pio_s1_arb_counter_enable) = '1' then 
        cal_dac_code_pio_s1_arb_share_counter <= cal_dac_code_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cal_dac_code_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cal_dac_code_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((cal_dac_code_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_cal_dac_code_pio_s1)) OR ((end_xfer_arb_share_counter_term_cal_dac_code_pio_s1 AND NOT cal_dac_code_pio_s1_non_bursting_master_requests)))) = '1' then 
        cal_dac_code_pio_s1_slavearbiterlockenable <= cal_dac_code_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_15/out cal_dac_code_pio/s1 arbiterlock, which is an e_assign
  nios2_clock_15_out_arbiterlock <= cal_dac_code_pio_s1_slavearbiterlockenable AND nios2_clock_15_out_continuerequest;
  --cal_dac_code_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cal_dac_code_pio_s1_slavearbiterlockenable2 <= cal_dac_code_pio_s1_arb_share_counter_next_value;
  --nios2_clock_15/out cal_dac_code_pio/s1 arbiterlock2, which is an e_assign
  nios2_clock_15_out_arbiterlock2 <= cal_dac_code_pio_s1_slavearbiterlockenable2 AND nios2_clock_15_out_continuerequest;
  --cal_dac_code_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  cal_dac_code_pio_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_15_out_continuerequest continued request, which is an e_assign
  nios2_clock_15_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 <= internal_nios2_clock_15_out_requests_cal_dac_code_pio_s1;
  --cal_dac_code_pio_s1_writedata mux, which is an e_mux
  cal_dac_code_pio_s1_writedata <= nios2_clock_15_out_writedata (13 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_clock_15_out_granted_cal_dac_code_pio_s1 <= internal_nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1;
  --nios2_clock_15/out saved-grant cal_dac_code_pio/s1, which is an e_assign
  nios2_clock_15_out_saved_grant_cal_dac_code_pio_s1 <= internal_nios2_clock_15_out_requests_cal_dac_code_pio_s1;
  --allow new arb cycle for cal_dac_code_pio/s1, which is an e_assign
  cal_dac_code_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  cal_dac_code_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  cal_dac_code_pio_s1_master_qreq_vector <= std_logic'('1');
  --cal_dac_code_pio_s1_reset_n assignment, which is an e_assign
  cal_dac_code_pio_s1_reset_n <= reset_n;
  cal_dac_code_pio_s1_chipselect <= internal_nios2_clock_15_out_granted_cal_dac_code_pio_s1;
  --cal_dac_code_pio_s1_firsttransfer first transaction, which is an e_assign
  cal_dac_code_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(cal_dac_code_pio_s1_begins_xfer) = '1'), cal_dac_code_pio_s1_unreg_firsttransfer, cal_dac_code_pio_s1_reg_firsttransfer);
  --cal_dac_code_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  cal_dac_code_pio_s1_unreg_firsttransfer <= NOT ((cal_dac_code_pio_s1_slavearbiterlockenable AND cal_dac_code_pio_s1_any_continuerequest));
  --cal_dac_code_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cal_dac_code_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cal_dac_code_pio_s1_begins_xfer) = '1' then 
        cal_dac_code_pio_s1_reg_firsttransfer <= cal_dac_code_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cal_dac_code_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cal_dac_code_pio_s1_beginbursttransfer_internal <= cal_dac_code_pio_s1_begins_xfer;
  --~cal_dac_code_pio_s1_write_n assignment, which is an e_mux
  cal_dac_code_pio_s1_write_n <= NOT ((internal_nios2_clock_15_out_granted_cal_dac_code_pio_s1 AND nios2_clock_15_out_write));
  --cal_dac_code_pio_s1_address mux, which is an e_mux
  cal_dac_code_pio_s1_address <= nios2_clock_15_out_nativeaddress;
  --d1_cal_dac_code_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cal_dac_code_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cal_dac_code_pio_s1_end_xfer <= cal_dac_code_pio_s1_end_xfer;
    end if;

  end process;

  --cal_dac_code_pio_s1_waits_for_read in a cycle, which is an e_mux
  cal_dac_code_pio_s1_waits_for_read <= cal_dac_code_pio_s1_in_a_read_cycle AND cal_dac_code_pio_s1_begins_xfer;
  --cal_dac_code_pio_s1_in_a_read_cycle assignment, which is an e_assign
  cal_dac_code_pio_s1_in_a_read_cycle <= internal_nios2_clock_15_out_granted_cal_dac_code_pio_s1 AND nios2_clock_15_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cal_dac_code_pio_s1_in_a_read_cycle;
  --cal_dac_code_pio_s1_waits_for_write in a cycle, which is an e_mux
  cal_dac_code_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cal_dac_code_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cal_dac_code_pio_s1_in_a_write_cycle assignment, which is an e_assign
  cal_dac_code_pio_s1_in_a_write_cycle <= internal_nios2_clock_15_out_granted_cal_dac_code_pio_s1 AND nios2_clock_15_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cal_dac_code_pio_s1_in_a_write_cycle;
  wait_for_cal_dac_code_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_15_out_granted_cal_dac_code_pio_s1 <= internal_nios2_clock_15_out_granted_cal_dac_code_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 <= internal_nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_15_out_requests_cal_dac_code_pio_s1 <= internal_nios2_clock_15_out_requests_cal_dac_code_pio_s1;
--synthesis translate_off
    --cal_dac_code_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity comparator_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal comparator_pio_s1_readdata : IN STD_LOGIC;
                 signal nios2_clock_11_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_11_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_11_out_read : IN STD_LOGIC;
                 signal nios2_clock_11_out_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal comparator_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal comparator_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal comparator_pio_s1_reset_n : OUT STD_LOGIC;
                 signal d1_comparator_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_11_out_granted_comparator_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_11_out_qualified_request_comparator_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_11_out_read_data_valid_comparator_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_11_out_requests_comparator_pio_s1 : OUT STD_LOGIC
              );
end entity comparator_pio_s1_arbitrator;


architecture europa of comparator_pio_s1_arbitrator is
                signal comparator_pio_s1_allgrants :  STD_LOGIC;
                signal comparator_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal comparator_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal comparator_pio_s1_any_continuerequest :  STD_LOGIC;
                signal comparator_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal comparator_pio_s1_arb_share_counter :  STD_LOGIC;
                signal comparator_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal comparator_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal comparator_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal comparator_pio_s1_begins_xfer :  STD_LOGIC;
                signal comparator_pio_s1_end_xfer :  STD_LOGIC;
                signal comparator_pio_s1_firsttransfer :  STD_LOGIC;
                signal comparator_pio_s1_grant_vector :  STD_LOGIC;
                signal comparator_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal comparator_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal comparator_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal comparator_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal comparator_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal comparator_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal comparator_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal comparator_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal comparator_pio_s1_waits_for_read :  STD_LOGIC;
                signal comparator_pio_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_comparator_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_11_out_granted_comparator_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_11_out_qualified_request_comparator_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_11_out_requests_comparator_pio_s1 :  STD_LOGIC;
                signal nios2_clock_11_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_11_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_11_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_11_out_saved_grant_comparator_pio_s1 :  STD_LOGIC;
                signal wait_for_comparator_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT comparator_pio_s1_end_xfer;
    end if;

  end process;

  comparator_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_11_out_qualified_request_comparator_pio_s1);
  --assign comparator_pio_s1_readdata_from_sa = comparator_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  comparator_pio_s1_readdata_from_sa <= comparator_pio_s1_readdata;
  internal_nios2_clock_11_out_requests_comparator_pio_s1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_11_out_read OR nios2_clock_11_out_write))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_11_out_read)))));
  --comparator_pio_s1_arb_share_counter set values, which is an e_mux
  comparator_pio_s1_arb_share_set_values <= std_logic'('1');
  --comparator_pio_s1_non_bursting_master_requests mux, which is an e_mux
  comparator_pio_s1_non_bursting_master_requests <= internal_nios2_clock_11_out_requests_comparator_pio_s1;
  --comparator_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  comparator_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --comparator_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  comparator_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(comparator_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(comparator_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(comparator_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(comparator_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --comparator_pio_s1_allgrants all slave grants, which is an e_mux
  comparator_pio_s1_allgrants <= comparator_pio_s1_grant_vector;
  --comparator_pio_s1_end_xfer assignment, which is an e_assign
  comparator_pio_s1_end_xfer <= NOT ((comparator_pio_s1_waits_for_read OR comparator_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_comparator_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_comparator_pio_s1 <= comparator_pio_s1_end_xfer AND (((NOT comparator_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --comparator_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  comparator_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_comparator_pio_s1 AND comparator_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_comparator_pio_s1 AND NOT comparator_pio_s1_non_bursting_master_requests));
  --comparator_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      comparator_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(comparator_pio_s1_arb_counter_enable) = '1' then 
        comparator_pio_s1_arb_share_counter <= comparator_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --comparator_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      comparator_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((comparator_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_comparator_pio_s1)) OR ((end_xfer_arb_share_counter_term_comparator_pio_s1 AND NOT comparator_pio_s1_non_bursting_master_requests)))) = '1' then 
        comparator_pio_s1_slavearbiterlockenable <= comparator_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_11/out comparator_pio/s1 arbiterlock, which is an e_assign
  nios2_clock_11_out_arbiterlock <= comparator_pio_s1_slavearbiterlockenable AND nios2_clock_11_out_continuerequest;
  --comparator_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  comparator_pio_s1_slavearbiterlockenable2 <= comparator_pio_s1_arb_share_counter_next_value;
  --nios2_clock_11/out comparator_pio/s1 arbiterlock2, which is an e_assign
  nios2_clock_11_out_arbiterlock2 <= comparator_pio_s1_slavearbiterlockenable2 AND nios2_clock_11_out_continuerequest;
  --comparator_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  comparator_pio_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_11_out_continuerequest continued request, which is an e_assign
  nios2_clock_11_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_11_out_qualified_request_comparator_pio_s1 <= internal_nios2_clock_11_out_requests_comparator_pio_s1;
  --master is always granted when requested
  internal_nios2_clock_11_out_granted_comparator_pio_s1 <= internal_nios2_clock_11_out_qualified_request_comparator_pio_s1;
  --nios2_clock_11/out saved-grant comparator_pio/s1, which is an e_assign
  nios2_clock_11_out_saved_grant_comparator_pio_s1 <= internal_nios2_clock_11_out_requests_comparator_pio_s1;
  --allow new arb cycle for comparator_pio/s1, which is an e_assign
  comparator_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  comparator_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  comparator_pio_s1_master_qreq_vector <= std_logic'('1');
  --comparator_pio_s1_reset_n assignment, which is an e_assign
  comparator_pio_s1_reset_n <= reset_n;
  --comparator_pio_s1_firsttransfer first transaction, which is an e_assign
  comparator_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(comparator_pio_s1_begins_xfer) = '1'), comparator_pio_s1_unreg_firsttransfer, comparator_pio_s1_reg_firsttransfer);
  --comparator_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  comparator_pio_s1_unreg_firsttransfer <= NOT ((comparator_pio_s1_slavearbiterlockenable AND comparator_pio_s1_any_continuerequest));
  --comparator_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      comparator_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(comparator_pio_s1_begins_xfer) = '1' then 
        comparator_pio_s1_reg_firsttransfer <= comparator_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --comparator_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  comparator_pio_s1_beginbursttransfer_internal <= comparator_pio_s1_begins_xfer;
  --comparator_pio_s1_address mux, which is an e_mux
  comparator_pio_s1_address <= nios2_clock_11_out_nativeaddress;
  --d1_comparator_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_comparator_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_comparator_pio_s1_end_xfer <= comparator_pio_s1_end_xfer;
    end if;

  end process;

  --comparator_pio_s1_waits_for_read in a cycle, which is an e_mux
  comparator_pio_s1_waits_for_read <= comparator_pio_s1_in_a_read_cycle AND comparator_pio_s1_begins_xfer;
  --comparator_pio_s1_in_a_read_cycle assignment, which is an e_assign
  comparator_pio_s1_in_a_read_cycle <= internal_nios2_clock_11_out_granted_comparator_pio_s1 AND nios2_clock_11_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= comparator_pio_s1_in_a_read_cycle;
  --comparator_pio_s1_waits_for_write in a cycle, which is an e_mux
  comparator_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(comparator_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --comparator_pio_s1_in_a_write_cycle assignment, which is an e_assign
  comparator_pio_s1_in_a_write_cycle <= internal_nios2_clock_11_out_granted_comparator_pio_s1 AND nios2_clock_11_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= comparator_pio_s1_in_a_write_cycle;
  wait_for_comparator_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_11_out_granted_comparator_pio_s1 <= internal_nios2_clock_11_out_granted_comparator_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_11_out_qualified_request_comparator_pio_s1 <= internal_nios2_clock_11_out_qualified_request_comparator_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_11_out_requests_comparator_pio_s1 <= internal_nios2_clock_11_out_requests_comparator_pio_s1;
--synthesis translate_off
    --comparator_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_0_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal cpu_0_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_reset_n : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_write : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_0_jtag_debug_module_end_xfer : OUT STD_LOGIC
              );
end entity cpu_0_jtag_debug_module_arbitrator;


architecture europa of cpu_0_jtag_debug_module_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_allgrants :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_0_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_cpu_0_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpu_0_jtag_debug_module_end_xfer;
    end if;

  end process;

  cpu_0_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module));
  --assign cpu_0_jtag_debug_module_readdata_from_sa = cpu_0_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_0_jtag_debug_module_readdata_from_sa <= cpu_0_jtag_debug_module_readdata;
  internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1000000010000100000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --cpu_0_jtag_debug_module_arb_share_counter set values, which is an e_mux
  cpu_0_jtag_debug_module_arb_share_set_values <= std_logic_vector'("01");
  --cpu_0_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  cpu_0_jtag_debug_module_non_bursting_master_requests <= ((internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module OR internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module) OR internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module) OR internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  --cpu_0_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  cpu_0_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --cpu_0_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  cpu_0_jtag_debug_module_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(cpu_0_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (cpu_0_jtag_debug_module_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(cpu_0_jtag_debug_module_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (cpu_0_jtag_debug_module_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --cpu_0_jtag_debug_module_allgrants all slave grants, which is an e_mux
  cpu_0_jtag_debug_module_allgrants <= (((or_reduce(cpu_0_jtag_debug_module_grant_vector)) OR (or_reduce(cpu_0_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_0_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_0_jtag_debug_module_grant_vector));
  --cpu_0_jtag_debug_module_end_xfer assignment, which is an e_assign
  cpu_0_jtag_debug_module_end_xfer <= NOT ((cpu_0_jtag_debug_module_waits_for_read OR cpu_0_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_end_xfer AND (((NOT cpu_0_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpu_0_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  cpu_0_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module AND cpu_0_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module AND NOT cpu_0_jtag_debug_module_non_bursting_master_requests));
  --cpu_0_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_0_jtag_debug_module_arb_counter_enable) = '1' then 
        cpu_0_jtag_debug_module_arb_share_counter <= cpu_0_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(cpu_0_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module AND NOT cpu_0_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        cpu_0_jtag_debug_module_slavearbiterlockenable <= or_reduce(cpu_0_jtag_debug_module_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= cpu_0_jtag_debug_module_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --cpu_0_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpu_0_jtag_debug_module_slavearbiterlockenable2 <= or_reduce(cpu_0_jtag_debug_module_arb_share_counter_next_value);
  --cpu_0/data_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= cpu_0_jtag_debug_module_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= cpu_0_jtag_debug_module_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= cpu_0_jtag_debug_module_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master granted cpu_0/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_0_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module))))));
    end if;

  end process;

  --cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  cpu_0_instruction_master_continuerequest <= last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module AND internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  --cpu_0_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  cpu_0_jtag_debug_module_any_continuerequest <= cpu_0_instruction_master_continuerequest OR cpu_0_data_master_continuerequest;
  internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module AND NOT ((((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR cpu_0_instruction_master_arbiterlock));
  --local readdatavalid cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module, which is an e_mux
  cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module <= (internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module AND cpu_0_data_master_read) AND NOT cpu_0_jtag_debug_module_waits_for_read;
  --cpu_0_jtag_debug_module_writedata mux, which is an e_mux
  cpu_0_jtag_debug_module_writedata <= cpu_0_data_master_writedata;
  internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(24 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1000000010000100000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --cpu_0/data_master granted cpu_0/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_0_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module))))));
    end if;

  end process;

  --cpu_0_data_master_continuerequest continued request, which is an e_mux
  cpu_0_data_master_continuerequest <= last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module AND internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module AND NOT ((((cpu_0_instruction_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR cpu_0_data_master_arbiterlock));
  --local readdatavalid cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module, which is an e_mux
  cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module <= (internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module AND cpu_0_instruction_master_read) AND NOT cpu_0_jtag_debug_module_waits_for_read;
  --allow new arb cycle for cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_jtag_debug_module_allow_new_arb_cycle <= NOT cpu_0_data_master_arbiterlock AND NOT cpu_0_instruction_master_arbiterlock;
  --cpu_0/instruction_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_jtag_debug_module_master_qreq_vector(0) <= internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  --cpu_0/instruction_master grant cpu_0/jtag_debug_module, which is an e_assign
  internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_grant_vector(0);
  --cpu_0/instruction_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_arb_winner(0) AND internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  --cpu_0/data_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_jtag_debug_module_master_qreq_vector(1) <= internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  --cpu_0/data_master grant cpu_0/jtag_debug_module, which is an e_assign
  internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_grant_vector(1);
  --cpu_0/data_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_arb_winner(1) AND internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  --cpu_0/jtag_debug_module chosen-master double-vector, which is an e_assign
  cpu_0_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((cpu_0_jtag_debug_module_master_qreq_vector & cpu_0_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT cpu_0_jtag_debug_module_master_qreq_vector & NOT cpu_0_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (cpu_0_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  cpu_0_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((cpu_0_jtag_debug_module_allow_new_arb_cycle AND or_reduce(cpu_0_jtag_debug_module_grant_vector)))) = '1'), cpu_0_jtag_debug_module_grant_vector, cpu_0_jtag_debug_module_saved_chosen_master_vector);
  --saved cpu_0_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_0_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        cpu_0_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(cpu_0_jtag_debug_module_grant_vector)) = '1'), cpu_0_jtag_debug_module_grant_vector, cpu_0_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  cpu_0_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((cpu_0_jtag_debug_module_chosen_master_double_vector(1) OR cpu_0_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((cpu_0_jtag_debug_module_chosen_master_double_vector(0) OR cpu_0_jtag_debug_module_chosen_master_double_vector(2)))));
  --cpu_0/jtag_debug_module chosen master rotated left, which is an e_assign
  cpu_0_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(cpu_0_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(cpu_0_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --cpu_0/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(cpu_0_jtag_debug_module_grant_vector)) = '1' then 
        cpu_0_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(cpu_0_jtag_debug_module_end_xfer) = '1'), cpu_0_jtag_debug_module_chosen_master_rot_left, cpu_0_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  cpu_0_jtag_debug_module_begintransfer <= cpu_0_jtag_debug_module_begins_xfer;
  --cpu_0_jtag_debug_module_reset_n assignment, which is an e_assign
  cpu_0_jtag_debug_module_reset_n <= reset_n;
  --assign cpu_0_jtag_debug_module_resetrequest_from_sa = cpu_0_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_0_jtag_debug_module_resetrequest_from_sa <= cpu_0_jtag_debug_module_resetrequest;
  cpu_0_jtag_debug_module_chipselect <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module OR internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  --cpu_0_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  cpu_0_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(cpu_0_jtag_debug_module_begins_xfer) = '1'), cpu_0_jtag_debug_module_unreg_firsttransfer, cpu_0_jtag_debug_module_reg_firsttransfer);
  --cpu_0_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  cpu_0_jtag_debug_module_unreg_firsttransfer <= NOT ((cpu_0_jtag_debug_module_slavearbiterlockenable AND cpu_0_jtag_debug_module_any_continuerequest));
  --cpu_0_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_0_jtag_debug_module_begins_xfer) = '1' then 
        cpu_0_jtag_debug_module_reg_firsttransfer <= cpu_0_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpu_0_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpu_0_jtag_debug_module_beginbursttransfer_internal <= cpu_0_jtag_debug_module_begins_xfer;
  --cpu_0_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  cpu_0_jtag_debug_module_arbitration_holdoff_internal <= cpu_0_jtag_debug_module_begins_xfer AND cpu_0_jtag_debug_module_firsttransfer;
  --cpu_0_jtag_debug_module_write assignment, which is an e_mux
  cpu_0_jtag_debug_module_write <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module AND cpu_0_data_master_write;
  shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --cpu_0_jtag_debug_module_address mux, which is an e_mux
  cpu_0_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master <= cpu_0_instruction_master_address_to_slave;
  --d1_cpu_0_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpu_0_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpu_0_jtag_debug_module_end_xfer <= cpu_0_jtag_debug_module_end_xfer;
    end if;

  end process;

  --cpu_0_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  cpu_0_jtag_debug_module_waits_for_read <= cpu_0_jtag_debug_module_in_a_read_cycle AND cpu_0_jtag_debug_module_begins_xfer;
  --cpu_0_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  cpu_0_jtag_debug_module_in_a_read_cycle <= ((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module AND cpu_0_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpu_0_jtag_debug_module_in_a_read_cycle;
  --cpu_0_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  cpu_0_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cpu_0_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  cpu_0_jtag_debug_module_in_a_write_cycle <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpu_0_jtag_debug_module_in_a_write_cycle;
  wait_for_cpu_0_jtag_debug_module_counter <= std_logic'('0');
  --cpu_0_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  cpu_0_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  cpu_0_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
--synthesis translate_off
    --cpu_0/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module;


architecture europa of jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module;


architecture europa of sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_0_data_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_byteenable_nios2_clock_9_in : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_10_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_11_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_12_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_13_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_14_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_15_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_16_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_17_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_18_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_2_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_3_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_4_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_5_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_6_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_7_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_nios2_clock_9_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_10_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_11_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_12_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_13_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_14_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_15_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_16_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_17_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_18_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_2_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_3_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_4_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_5_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_6_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_7_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_9_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_10_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_11_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_12_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_13_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_14_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_15_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_16_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_17_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_18_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_2_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_3_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_4_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_5_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_6_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_7_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_9_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_10_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_11_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_12_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_13_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_14_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_15_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_16_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_17_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_18_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_2_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_3_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_4_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_5_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_6_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_7_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_9_in : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_10_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_11_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_12_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_13_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_14_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_15_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_16_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_17_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_18_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_1_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_2_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_3_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_4_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_5_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_6_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_7_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_9_in_end_xfer : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal nios2_clock_10_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_10_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_11_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_11_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_12_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_12_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_13_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_13_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_14_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_14_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_15_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_15_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_16_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_16_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_17_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_17_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_18_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_18_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_2_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_2_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_3_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_3_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_4_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_4_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_5_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_5_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_6_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_6_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_7_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_7_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_9_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_9_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal processor_clk : IN STD_LOGIC;
                 signal processor_clk_reset_n : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_0_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_0_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : OUT STD_LOGIC;
                 signal cpu_0_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_data_master_readdatavalid : OUT STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_0_data_master_arbitrator;


architecture europa of cpu_0_data_master_arbitrator is
component jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module;

component sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module;

                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_0_data_master_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_0_data_master_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_0_data_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_data_master_is_granted_some_slave :  STD_LOGIC;
                signal cpu_0_data_master_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_0_data_master_read_last_time :  STD_LOGIC;
                signal cpu_0_data_master_run :  STD_LOGIC;
                signal cpu_0_data_master_write_last_time :  STD_LOGIC;
                signal cpu_0_data_master_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal internal_cpu_0_data_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_cpu_0_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_0_data_master_latency_counter :  STD_LOGIC;
                signal internal_cpu_0_data_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_cpu_0_data_master_latency_counter :  STD_LOGIC;
                signal p1_dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_cpu_0_data_master_readdatavalid :  STD_LOGIC;
                signal processor_clk_jtag_uart_0_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal processor_clk_sys_clk_timer_s1_irq_from_sa :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_requests_cpu_0_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_granted_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpu_0_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_1_in OR NOT cpu_0_data_master_requests_nios2_clock_1_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_1_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_1_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_10_in OR NOT cpu_0_data_master_requests_nios2_clock_10_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_10_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_10_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_10_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_10_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_11_in OR NOT cpu_0_data_master_requests_nios2_clock_11_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_11_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_11_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_11_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_11_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_12_in OR NOT cpu_0_data_master_requests_nios2_clock_12_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_12_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_12_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_0_data_master_run <= ((r_0 AND r_1) AND r_2) AND r_3;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_12_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_12_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_13_in OR NOT cpu_0_data_master_requests_nios2_clock_13_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_13_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_13_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_13_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_13_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_14_in OR NOT cpu_0_data_master_requests_nios2_clock_14_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_14_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_14_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_14_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_14_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_15_in OR NOT cpu_0_data_master_requests_nios2_clock_15_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_15_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_15_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_15_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_15_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_16_in OR NOT cpu_0_data_master_requests_nios2_clock_16_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_16_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_16_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_16_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_16_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_17_in OR NOT cpu_0_data_master_requests_nios2_clock_17_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_17_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_17_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_17_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_17_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_18_in OR NOT cpu_0_data_master_requests_nios2_clock_18_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_18_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_18_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_18_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_18_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_2_in OR NOT cpu_0_data_master_requests_nios2_clock_2_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_2_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_2_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_2_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_2_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_3_in OR NOT cpu_0_data_master_requests_nios2_clock_3_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_3_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_3_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_3_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_3_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_4_in OR NOT cpu_0_data_master_requests_nios2_clock_4_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_4_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_4_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_4_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_4_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_5_in OR NOT cpu_0_data_master_requests_nios2_clock_5_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_5_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_5_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))));
  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_5_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_5_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_6_in OR NOT cpu_0_data_master_requests_nios2_clock_6_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_6_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_6_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_6_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_6_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_nios2_clock_7_in OR NOT cpu_0_data_master_requests_nios2_clock_7_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_7_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_7_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_7_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_7_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_data_master_qualified_request_nios2_clock_9_in OR (((cpu_0_data_master_write AND NOT(or_reduce(cpu_0_data_master_byteenable_nios2_clock_9_in))) AND internal_cpu_0_data_master_dbs_address(1)))) OR NOT cpu_0_data_master_requests_nios2_clock_9_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_9_in OR NOT cpu_0_data_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_9_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_0_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_nios2_clock_9_in OR NOT cpu_0_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_9_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_0_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_write)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_0_data_master_address_to_slave <= cpu_0_data_master_address(24 DOWNTO 0);
  --cpu_0_data_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_data_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_0_data_master_read_but_no_slave_selected <= (cpu_0_data_master_read AND cpu_0_data_master_run) AND NOT cpu_0_data_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_0_data_master_is_granted_some_slave <= ((((((((((((((((cpu_0_data_master_granted_cpu_0_jtag_debug_module OR cpu_0_data_master_granted_nios2_clock_1_in) OR cpu_0_data_master_granted_nios2_clock_10_in) OR cpu_0_data_master_granted_nios2_clock_11_in) OR cpu_0_data_master_granted_nios2_clock_12_in) OR cpu_0_data_master_granted_nios2_clock_13_in) OR cpu_0_data_master_granted_nios2_clock_14_in) OR cpu_0_data_master_granted_nios2_clock_15_in) OR cpu_0_data_master_granted_nios2_clock_16_in) OR cpu_0_data_master_granted_nios2_clock_17_in) OR cpu_0_data_master_granted_nios2_clock_18_in) OR cpu_0_data_master_granted_nios2_clock_2_in) OR cpu_0_data_master_granted_nios2_clock_3_in) OR cpu_0_data_master_granted_nios2_clock_4_in) OR cpu_0_data_master_granted_nios2_clock_5_in) OR cpu_0_data_master_granted_nios2_clock_6_in) OR cpu_0_data_master_granted_nios2_clock_7_in) OR cpu_0_data_master_granted_nios2_clock_9_in;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_0_data_master_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_0_data_master_readdatavalid <= ((((((((((((((((((((((((((((((((((((((((((((((((((((cpu_0_data_master_read_but_no_slave_selected OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_1_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_10_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_11_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_12_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_13_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_14_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_15_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_16_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_17_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_18_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_2_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_3_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_4_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_5_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_6_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR cpu_0_data_master_read_data_valid_nios2_clock_7_in) OR cpu_0_data_master_read_but_no_slave_selected) OR pre_flush_cpu_0_data_master_readdatavalid) OR ((cpu_0_data_master_read_data_valid_nios2_clock_9_in AND dbs_counter_overflow));
  --cpu_0/data_master readdata mux, which is an e_mux
  cpu_0_data_master_readdata <= ((((((((((((((((((A_REP(NOT ((cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module AND cpu_0_data_master_read)) , 32) OR cpu_0_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_1_in AND cpu_0_data_master_read)) , 32) OR nios2_clock_1_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_10_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (nios2_clock_10_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_11_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (nios2_clock_11_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_12_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (nios2_clock_12_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_13_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (nios2_clock_13_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_14_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (nios2_clock_14_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_15_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("0000000000000000") & (nios2_clock_15_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_16_in AND cpu_0_data_master_read)) , 32) OR nios2_clock_16_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_17_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (nios2_clock_17_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_18_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (nios2_clock_18_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_2_in AND cpu_0_data_master_read)) , 32) OR nios2_clock_2_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_3_in AND cpu_0_data_master_read)) , 32) OR (std_logic_vector'("0000000000000000") & (nios2_clock_3_in_readdata_from_sa))))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_4_in AND cpu_0_data_master_read)) , 32) OR nios2_clock_4_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_5_in AND cpu_0_data_master_read)) , 32) OR nios2_clock_5_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_6_in AND cpu_0_data_master_read)) , 32) OR nios2_clock_6_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_7_in AND cpu_0_data_master_read)) , 32) OR nios2_clock_7_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_data_master_qualified_request_nios2_clock_9_in AND cpu_0_data_master_read)) , 32) OR Std_Logic_Vector'(nios2_clock_9_in_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0)));
  --actual waitrequest port, which is an e_assign
  internal_cpu_0_data_master_waitrequest <= NOT cpu_0_data_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_0_data_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_cpu_0_data_master_latency_counter <= p1_cpu_0_data_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_0_data_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((cpu_0_data_master_run AND cpu_0_data_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_cpu_0_data_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --jtag_uart_0_avalon_jtag_slave_irq_from_sa from altpll_0_c0 to processor_clk
  jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master : jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module
    port map(
      data_out => processor_clk_jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      clk => processor_clk,
      data_in => jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      reset_n => processor_clk_reset_n
    );


  --irq assign, which is an e_assign
  cpu_0_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(processor_clk_sys_clk_timer_s1_irq_from_sa) & A_ToStdLogicVector(processor_clk_jtag_uart_0_avalon_jtag_slave_irq_from_sa));
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((((((NOT std_logic_vector'("00000000000000000000000000000000")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_requests_nios2_clock_9_in)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_write)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT(or_reduce(cpu_0_data_master_byteenable_nios2_clock_9_in))))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_0_data_master_granted_nios2_clock_9_in AND cpu_0_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_9_in_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_0_data_master_granted_nios2_clock_9_in AND cpu_0_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_9_in_waitrequest_from_sa)))))));
  --input to dbs-16 stored 0, which is an e_mux
  p1_dbs_16_reg_segment_0 <= nios2_clock_9_in_readdata_from_sa;
  --dbs register for dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_0_data_master_dbs_address(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
      end if;
    end if;

  end process;

  --mux write dbs 1, which is an e_mux
  cpu_0_data_master_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_dbs_address(1))) = '1'), cpu_0_data_master_writedata(31 DOWNTO 16), cpu_0_data_master_writedata(15 DOWNTO 0));
  --dbs count increment, which is an e_mux
  cpu_0_data_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_0_data_master_requests_nios2_clock_9_in)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_cpu_0_data_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_cpu_0_data_master_dbs_address)) + (std_logic_vector'("0") & (cpu_0_data_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_0_data_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_cpu_0_data_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_irq_from_sa from clk_0 to processor_clk
  sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master : sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module
    port map(
      data_out => processor_clk_sys_clk_timer_s1_irq_from_sa,
      clk => processor_clk,
      data_in => sys_clk_timer_s1_irq_from_sa,
      reset_n => processor_clk_reset_n
    );


  --vhdl renameroo for output signals
  cpu_0_data_master_address_to_slave <= internal_cpu_0_data_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_0_data_master_dbs_address <= internal_cpu_0_data_master_dbs_address;
  --vhdl renameroo for output signals
  cpu_0_data_master_latency_counter <= internal_cpu_0_data_master_latency_counter;
  --vhdl renameroo for output signals
  cpu_0_data_master_waitrequest <= internal_cpu_0_data_master_waitrequest;
--synthesis translate_off
    --cpu_0_data_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_data_master_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_0_data_master_address_last_time <= cpu_0_data_master_address;
      end if;

    end process;

    --cpu_0/data_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_0_data_master_waitrequest AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
      end if;

    end process;

    --cpu_0_data_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_0_data_master_address /= cpu_0_data_master_address_last_time))))) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("cpu_0_data_master_address did not heed wait!!!"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_0_data_master_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_data_master_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        cpu_0_data_master_byteenable_last_time <= cpu_0_data_master_byteenable;
      end if;

    end process;

    --cpu_0_data_master_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_0_data_master_byteenable /= cpu_0_data_master_byteenable_last_time))))) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("cpu_0_data_master_byteenable did not heed wait!!!"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_0_data_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_data_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_0_data_master_read_last_time <= cpu_0_data_master_read;
      end if;

    end process;

    --cpu_0_data_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_0_data_master_read) /= std_logic'(cpu_0_data_master_read_last_time)))))) = '1' then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("cpu_0_data_master_read did not heed wait!!!"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_0_data_master_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_data_master_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_0_data_master_write_last_time <= cpu_0_data_master_write;
      end if;

    end process;

    --cpu_0_data_master_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_0_data_master_write) /= std_logic'(cpu_0_data_master_write_last_time)))))) = '1' then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("cpu_0_data_master_write did not heed wait!!!"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_0_data_master_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_data_master_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_0_data_master_writedata_last_time <= cpu_0_data_master_writedata;
      end if;

    end process;

    --cpu_0_data_master_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((cpu_0_data_master_writedata /= cpu_0_data_master_writedata_last_time)))) AND cpu_0_data_master_write)) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("cpu_0_data_master_writedata did not heed wait!!!"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_0_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_instruction_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_granted_nios2_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_instruction_master_granted_nios2_clock_8_in : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_nios2_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_nios2_clock_8_in : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_nios2_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_nios2_clock_8_in : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_nios2_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_nios2_clock_8_in : IN STD_LOGIC;
                 signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_0_in_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_clock_8_in_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_8_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_8_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_0_instruction_master_latency_counter : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_0_instruction_master_arbitrator;


architecture europa of cpu_0_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_0_instruction_master_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_0_instruction_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal cpu_0_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_0_instruction_master_read_last_time :  STD_LOGIC;
                signal cpu_0_instruction_master_run :  STD_LOGIC;
                signal dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_cpu_0_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_0_instruction_master_latency_counter :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_cpu_0_instruction_master_latency_counter :  STD_LOGIC;
                signal p1_dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_cpu_0_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_instruction_master_requests_cpu_0_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_granted_cpu_0_jtag_debug_module OR NOT cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpu_0_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_qualified_request_nios2_clock_0_in OR NOT cpu_0_instruction_master_requests_nios2_clock_0_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_instruction_master_qualified_request_nios2_clock_0_in OR NOT (cpu_0_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_0_instruction_master_read))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_0_instruction_master_run <= r_0 AND r_3;
  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_qualified_request_nios2_clock_8_in OR NOT cpu_0_instruction_master_requests_nios2_clock_8_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_instruction_master_qualified_request_nios2_clock_8_in OR NOT cpu_0_instruction_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_8_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_0_instruction_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_read)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_0_instruction_master_address_to_slave <= cpu_0_instruction_master_address(24 DOWNTO 0);
  --cpu_0_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_0_instruction_master_read_but_no_slave_selected <= (cpu_0_instruction_master_read AND cpu_0_instruction_master_run) AND NOT cpu_0_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_0_instruction_master_is_granted_some_slave <= (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module OR cpu_0_instruction_master_granted_nios2_clock_0_in) OR cpu_0_instruction_master_granted_nios2_clock_8_in;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_0_instruction_master_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_0_instruction_master_readdatavalid <= (((((((cpu_0_instruction_master_read_but_no_slave_selected OR pre_flush_cpu_0_instruction_master_readdatavalid) OR cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module) OR cpu_0_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_0_instruction_master_readdatavalid) OR cpu_0_instruction_master_read_data_valid_nios2_clock_0_in) OR cpu_0_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_0_instruction_master_readdatavalid) OR ((cpu_0_instruction_master_read_data_valid_nios2_clock_8_in AND dbs_counter_overflow));
  --cpu_0/instruction_master readdata mux, which is an e_mux
  cpu_0_instruction_master_readdata <= (((A_REP(NOT ((cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module AND cpu_0_instruction_master_read)) , 32) OR cpu_0_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT ((cpu_0_instruction_master_qualified_request_nios2_clock_0_in AND cpu_0_instruction_master_read)) , 32) OR nios2_clock_0_in_readdata_from_sa))) AND ((A_REP(NOT ((cpu_0_instruction_master_qualified_request_nios2_clock_8_in AND cpu_0_instruction_master_read)) , 32) OR Std_Logic_Vector'(nios2_clock_8_in_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0)));
  --actual waitrequest port, which is an e_assign
  internal_cpu_0_instruction_master_waitrequest <= NOT cpu_0_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_0_instruction_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_cpu_0_instruction_master_latency_counter <= p1_cpu_0_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_0_instruction_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((cpu_0_instruction_master_run AND cpu_0_instruction_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_cpu_0_instruction_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_cpu_0_instruction_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --input to dbs-16 stored 0, which is an e_mux
  p1_dbs_16_reg_segment_0 <= nios2_clock_8_in_readdata_from_sa;
  --dbs register for dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_0_instruction_master_dbs_address(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
      end if;
    end if;

  end process;

  --dbs count increment, which is an e_mux
  cpu_0_instruction_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_0_instruction_master_requests_nios2_clock_8_in)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_cpu_0_instruction_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_cpu_0_instruction_master_dbs_address)) + (std_logic_vector'("0") & (cpu_0_instruction_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_0_instruction_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_cpu_0_instruction_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_0_instruction_master_granted_nios2_clock_8_in AND cpu_0_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_clock_8_in_waitrequest_from_sa)))));
  --vhdl renameroo for output signals
  cpu_0_instruction_master_address_to_slave <= internal_cpu_0_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_dbs_address <= internal_cpu_0_instruction_master_dbs_address;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_latency_counter <= internal_cpu_0_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_waitrequest <= internal_cpu_0_instruction_master_waitrequest;
--synthesis translate_off
    --cpu_0_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_instruction_master_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_0_instruction_master_address_last_time <= cpu_0_instruction_master_address;
      end if;

    end process;

    --cpu_0/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_0_instruction_master_waitrequest AND (cpu_0_instruction_master_read);
      end if;

    end process;

    --cpu_0_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_0_instruction_master_address /= cpu_0_instruction_master_address_last_time))))) = '1' then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("cpu_0_instruction_master_address did not heed wait!!!"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_0_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_0_instruction_master_read_last_time <= cpu_0_instruction_master_read;
      end if;

    end process;

    --cpu_0_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_0_instruction_master_read) /= std_logic'(cpu_0_instruction_master_read_last_time)))))) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("cpu_0_instruction_master_read did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gen_code_strobe_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal gen_code_strobe_s1_readdata : IN STD_LOGIC;
                 signal nios2_clock_13_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_13_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_13_out_read : IN STD_LOGIC;
                 signal nios2_clock_13_out_write : IN STD_LOGIC;
                 signal nios2_clock_13_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_gen_code_strobe_s1_end_xfer : OUT STD_LOGIC;
                 signal gen_code_strobe_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gen_code_strobe_s1_chipselect : OUT STD_LOGIC;
                 signal gen_code_strobe_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal gen_code_strobe_s1_reset_n : OUT STD_LOGIC;
                 signal gen_code_strobe_s1_write_n : OUT STD_LOGIC;
                 signal gen_code_strobe_s1_writedata : OUT STD_LOGIC;
                 signal nios2_clock_13_out_granted_gen_code_strobe_s1 : OUT STD_LOGIC;
                 signal nios2_clock_13_out_qualified_request_gen_code_strobe_s1 : OUT STD_LOGIC;
                 signal nios2_clock_13_out_read_data_valid_gen_code_strobe_s1 : OUT STD_LOGIC;
                 signal nios2_clock_13_out_requests_gen_code_strobe_s1 : OUT STD_LOGIC
              );
end entity gen_code_strobe_s1_arbitrator;


architecture europa of gen_code_strobe_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gen_code_strobe_s1 :  STD_LOGIC;
                signal gen_code_strobe_s1_allgrants :  STD_LOGIC;
                signal gen_code_strobe_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal gen_code_strobe_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gen_code_strobe_s1_any_continuerequest :  STD_LOGIC;
                signal gen_code_strobe_s1_arb_counter_enable :  STD_LOGIC;
                signal gen_code_strobe_s1_arb_share_counter :  STD_LOGIC;
                signal gen_code_strobe_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal gen_code_strobe_s1_arb_share_set_values :  STD_LOGIC;
                signal gen_code_strobe_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal gen_code_strobe_s1_begins_xfer :  STD_LOGIC;
                signal gen_code_strobe_s1_end_xfer :  STD_LOGIC;
                signal gen_code_strobe_s1_firsttransfer :  STD_LOGIC;
                signal gen_code_strobe_s1_grant_vector :  STD_LOGIC;
                signal gen_code_strobe_s1_in_a_read_cycle :  STD_LOGIC;
                signal gen_code_strobe_s1_in_a_write_cycle :  STD_LOGIC;
                signal gen_code_strobe_s1_master_qreq_vector :  STD_LOGIC;
                signal gen_code_strobe_s1_non_bursting_master_requests :  STD_LOGIC;
                signal gen_code_strobe_s1_reg_firsttransfer :  STD_LOGIC;
                signal gen_code_strobe_s1_slavearbiterlockenable :  STD_LOGIC;
                signal gen_code_strobe_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal gen_code_strobe_s1_unreg_firsttransfer :  STD_LOGIC;
                signal gen_code_strobe_s1_waits_for_read :  STD_LOGIC;
                signal gen_code_strobe_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_13_out_granted_gen_code_strobe_s1 :  STD_LOGIC;
                signal internal_nios2_clock_13_out_qualified_request_gen_code_strobe_s1 :  STD_LOGIC;
                signal internal_nios2_clock_13_out_requests_gen_code_strobe_s1 :  STD_LOGIC;
                signal nios2_clock_13_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_13_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_13_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_13_out_saved_grant_gen_code_strobe_s1 :  STD_LOGIC;
                signal wait_for_gen_code_strobe_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gen_code_strobe_s1_end_xfer;
    end if;

  end process;

  gen_code_strobe_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_13_out_qualified_request_gen_code_strobe_s1);
  --assign gen_code_strobe_s1_readdata_from_sa = gen_code_strobe_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gen_code_strobe_s1_readdata_from_sa <= gen_code_strobe_s1_readdata;
  internal_nios2_clock_13_out_requests_gen_code_strobe_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_13_out_read OR nios2_clock_13_out_write)))))));
  --gen_code_strobe_s1_arb_share_counter set values, which is an e_mux
  gen_code_strobe_s1_arb_share_set_values <= std_logic'('1');
  --gen_code_strobe_s1_non_bursting_master_requests mux, which is an e_mux
  gen_code_strobe_s1_non_bursting_master_requests <= internal_nios2_clock_13_out_requests_gen_code_strobe_s1;
  --gen_code_strobe_s1_any_bursting_master_saved_grant mux, which is an e_mux
  gen_code_strobe_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --gen_code_strobe_s1_arb_share_counter_next_value assignment, which is an e_assign
  gen_code_strobe_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gen_code_strobe_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_strobe_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gen_code_strobe_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_strobe_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gen_code_strobe_s1_allgrants all slave grants, which is an e_mux
  gen_code_strobe_s1_allgrants <= gen_code_strobe_s1_grant_vector;
  --gen_code_strobe_s1_end_xfer assignment, which is an e_assign
  gen_code_strobe_s1_end_xfer <= NOT ((gen_code_strobe_s1_waits_for_read OR gen_code_strobe_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_gen_code_strobe_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gen_code_strobe_s1 <= gen_code_strobe_s1_end_xfer AND (((NOT gen_code_strobe_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gen_code_strobe_s1_arb_share_counter arbitration counter enable, which is an e_assign
  gen_code_strobe_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gen_code_strobe_s1 AND gen_code_strobe_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_gen_code_strobe_s1 AND NOT gen_code_strobe_s1_non_bursting_master_requests));
  --gen_code_strobe_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_strobe_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gen_code_strobe_s1_arb_counter_enable) = '1' then 
        gen_code_strobe_s1_arb_share_counter <= gen_code_strobe_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gen_code_strobe_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_strobe_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gen_code_strobe_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_gen_code_strobe_s1)) OR ((end_xfer_arb_share_counter_term_gen_code_strobe_s1 AND NOT gen_code_strobe_s1_non_bursting_master_requests)))) = '1' then 
        gen_code_strobe_s1_slavearbiterlockenable <= gen_code_strobe_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_13/out gen_code_strobe/s1 arbiterlock, which is an e_assign
  nios2_clock_13_out_arbiterlock <= gen_code_strobe_s1_slavearbiterlockenable AND nios2_clock_13_out_continuerequest;
  --gen_code_strobe_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gen_code_strobe_s1_slavearbiterlockenable2 <= gen_code_strobe_s1_arb_share_counter_next_value;
  --nios2_clock_13/out gen_code_strobe/s1 arbiterlock2, which is an e_assign
  nios2_clock_13_out_arbiterlock2 <= gen_code_strobe_s1_slavearbiterlockenable2 AND nios2_clock_13_out_continuerequest;
  --gen_code_strobe_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  gen_code_strobe_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_13_out_continuerequest continued request, which is an e_assign
  nios2_clock_13_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_13_out_qualified_request_gen_code_strobe_s1 <= internal_nios2_clock_13_out_requests_gen_code_strobe_s1;
  --gen_code_strobe_s1_writedata mux, which is an e_mux
  gen_code_strobe_s1_writedata <= nios2_clock_13_out_writedata(0);
  --master is always granted when requested
  internal_nios2_clock_13_out_granted_gen_code_strobe_s1 <= internal_nios2_clock_13_out_qualified_request_gen_code_strobe_s1;
  --nios2_clock_13/out saved-grant gen_code_strobe/s1, which is an e_assign
  nios2_clock_13_out_saved_grant_gen_code_strobe_s1 <= internal_nios2_clock_13_out_requests_gen_code_strobe_s1;
  --allow new arb cycle for gen_code_strobe/s1, which is an e_assign
  gen_code_strobe_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gen_code_strobe_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gen_code_strobe_s1_master_qreq_vector <= std_logic'('1');
  --gen_code_strobe_s1_reset_n assignment, which is an e_assign
  gen_code_strobe_s1_reset_n <= reset_n;
  gen_code_strobe_s1_chipselect <= internal_nios2_clock_13_out_granted_gen_code_strobe_s1;
  --gen_code_strobe_s1_firsttransfer first transaction, which is an e_assign
  gen_code_strobe_s1_firsttransfer <= A_WE_StdLogic((std_logic'(gen_code_strobe_s1_begins_xfer) = '1'), gen_code_strobe_s1_unreg_firsttransfer, gen_code_strobe_s1_reg_firsttransfer);
  --gen_code_strobe_s1_unreg_firsttransfer first transaction, which is an e_assign
  gen_code_strobe_s1_unreg_firsttransfer <= NOT ((gen_code_strobe_s1_slavearbiterlockenable AND gen_code_strobe_s1_any_continuerequest));
  --gen_code_strobe_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_strobe_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gen_code_strobe_s1_begins_xfer) = '1' then 
        gen_code_strobe_s1_reg_firsttransfer <= gen_code_strobe_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gen_code_strobe_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gen_code_strobe_s1_beginbursttransfer_internal <= gen_code_strobe_s1_begins_xfer;
  --~gen_code_strobe_s1_write_n assignment, which is an e_mux
  gen_code_strobe_s1_write_n <= NOT ((internal_nios2_clock_13_out_granted_gen_code_strobe_s1 AND nios2_clock_13_out_write));
  --gen_code_strobe_s1_address mux, which is an e_mux
  gen_code_strobe_s1_address <= nios2_clock_13_out_nativeaddress;
  --d1_gen_code_strobe_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gen_code_strobe_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gen_code_strobe_s1_end_xfer <= gen_code_strobe_s1_end_xfer;
    end if;

  end process;

  --gen_code_strobe_s1_waits_for_read in a cycle, which is an e_mux
  gen_code_strobe_s1_waits_for_read <= gen_code_strobe_s1_in_a_read_cycle AND gen_code_strobe_s1_begins_xfer;
  --gen_code_strobe_s1_in_a_read_cycle assignment, which is an e_assign
  gen_code_strobe_s1_in_a_read_cycle <= internal_nios2_clock_13_out_granted_gen_code_strobe_s1 AND nios2_clock_13_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gen_code_strobe_s1_in_a_read_cycle;
  --gen_code_strobe_s1_waits_for_write in a cycle, which is an e_mux
  gen_code_strobe_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_strobe_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --gen_code_strobe_s1_in_a_write_cycle assignment, which is an e_assign
  gen_code_strobe_s1_in_a_write_cycle <= internal_nios2_clock_13_out_granted_gen_code_strobe_s1 AND nios2_clock_13_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gen_code_strobe_s1_in_a_write_cycle;
  wait_for_gen_code_strobe_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_13_out_granted_gen_code_strobe_s1 <= internal_nios2_clock_13_out_granted_gen_code_strobe_s1;
  --vhdl renameroo for output signals
  nios2_clock_13_out_qualified_request_gen_code_strobe_s1 <= internal_nios2_clock_13_out_qualified_request_gen_code_strobe_s1;
  --vhdl renameroo for output signals
  nios2_clock_13_out_requests_gen_code_strobe_s1 <= internal_nios2_clock_13_out_requests_gen_code_strobe_s1;
--synthesis translate_off
    --gen_code_strobe/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gen_code_value_pio_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal gen_code_value_pio_0_s1_readdata : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal nios2_clock_6_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_6_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_6_out_read : IN STD_LOGIC;
                 signal nios2_clock_6_out_write : IN STD_LOGIC;
                 signal nios2_clock_6_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_gen_code_value_pio_0_s1_end_xfer : OUT STD_LOGIC;
                 signal gen_code_value_pio_0_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gen_code_value_pio_0_s1_chipselect : OUT STD_LOGIC;
                 signal gen_code_value_pio_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal gen_code_value_pio_0_s1_reset_n : OUT STD_LOGIC;
                 signal gen_code_value_pio_0_s1_write_n : OUT STD_LOGIC;
                 signal gen_code_value_pio_0_s1_writedata : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal nios2_clock_6_out_granted_gen_code_value_pio_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_6_out_requests_gen_code_value_pio_0_s1 : OUT STD_LOGIC
              );
end entity gen_code_value_pio_0_s1_arbitrator;


architecture europa of gen_code_value_pio_0_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_allgrants :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_any_continuerequest :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_arb_counter_enable :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_arb_share_counter :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_arb_share_set_values :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_begins_xfer :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_end_xfer :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_firsttransfer :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_grant_vector :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_master_qreq_vector :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_waits_for_read :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_6_out_granted_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal internal_nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal internal_nios2_clock_6_out_requests_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal nios2_clock_6_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_6_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_6_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_6_out_saved_grant_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal wait_for_gen_code_value_pio_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gen_code_value_pio_0_s1_end_xfer;
    end if;

  end process;

  gen_code_value_pio_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1);
  --assign gen_code_value_pio_0_s1_readdata_from_sa = gen_code_value_pio_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gen_code_value_pio_0_s1_readdata_from_sa <= gen_code_value_pio_0_s1_readdata;
  internal_nios2_clock_6_out_requests_gen_code_value_pio_0_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_6_out_read OR nios2_clock_6_out_write)))))));
  --gen_code_value_pio_0_s1_arb_share_counter set values, which is an e_mux
  gen_code_value_pio_0_s1_arb_share_set_values <= std_logic'('1');
  --gen_code_value_pio_0_s1_non_bursting_master_requests mux, which is an e_mux
  gen_code_value_pio_0_s1_non_bursting_master_requests <= internal_nios2_clock_6_out_requests_gen_code_value_pio_0_s1;
  --gen_code_value_pio_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  gen_code_value_pio_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --gen_code_value_pio_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  gen_code_value_pio_0_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gen_code_value_pio_0_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_value_pio_0_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gen_code_value_pio_0_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_value_pio_0_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gen_code_value_pio_0_s1_allgrants all slave grants, which is an e_mux
  gen_code_value_pio_0_s1_allgrants <= gen_code_value_pio_0_s1_grant_vector;
  --gen_code_value_pio_0_s1_end_xfer assignment, which is an e_assign
  gen_code_value_pio_0_s1_end_xfer <= NOT ((gen_code_value_pio_0_s1_waits_for_read OR gen_code_value_pio_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_gen_code_value_pio_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gen_code_value_pio_0_s1 <= gen_code_value_pio_0_s1_end_xfer AND (((NOT gen_code_value_pio_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gen_code_value_pio_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  gen_code_value_pio_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gen_code_value_pio_0_s1 AND gen_code_value_pio_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_gen_code_value_pio_0_s1 AND NOT gen_code_value_pio_0_s1_non_bursting_master_requests));
  --gen_code_value_pio_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_value_pio_0_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gen_code_value_pio_0_s1_arb_counter_enable) = '1' then 
        gen_code_value_pio_0_s1_arb_share_counter <= gen_code_value_pio_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gen_code_value_pio_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_value_pio_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gen_code_value_pio_0_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_gen_code_value_pio_0_s1)) OR ((end_xfer_arb_share_counter_term_gen_code_value_pio_0_s1 AND NOT gen_code_value_pio_0_s1_non_bursting_master_requests)))) = '1' then 
        gen_code_value_pio_0_s1_slavearbiterlockenable <= gen_code_value_pio_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_6/out gen_code_value_pio_0/s1 arbiterlock, which is an e_assign
  nios2_clock_6_out_arbiterlock <= gen_code_value_pio_0_s1_slavearbiterlockenable AND nios2_clock_6_out_continuerequest;
  --gen_code_value_pio_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gen_code_value_pio_0_s1_slavearbiterlockenable2 <= gen_code_value_pio_0_s1_arb_share_counter_next_value;
  --nios2_clock_6/out gen_code_value_pio_0/s1 arbiterlock2, which is an e_assign
  nios2_clock_6_out_arbiterlock2 <= gen_code_value_pio_0_s1_slavearbiterlockenable2 AND nios2_clock_6_out_continuerequest;
  --gen_code_value_pio_0_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  gen_code_value_pio_0_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_6_out_continuerequest continued request, which is an e_assign
  nios2_clock_6_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 <= internal_nios2_clock_6_out_requests_gen_code_value_pio_0_s1;
  --gen_code_value_pio_0_s1_writedata mux, which is an e_mux
  gen_code_value_pio_0_s1_writedata <= nios2_clock_6_out_writedata (23 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_clock_6_out_granted_gen_code_value_pio_0_s1 <= internal_nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1;
  --nios2_clock_6/out saved-grant gen_code_value_pio_0/s1, which is an e_assign
  nios2_clock_6_out_saved_grant_gen_code_value_pio_0_s1 <= internal_nios2_clock_6_out_requests_gen_code_value_pio_0_s1;
  --allow new arb cycle for gen_code_value_pio_0/s1, which is an e_assign
  gen_code_value_pio_0_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gen_code_value_pio_0_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gen_code_value_pio_0_s1_master_qreq_vector <= std_logic'('1');
  --gen_code_value_pio_0_s1_reset_n assignment, which is an e_assign
  gen_code_value_pio_0_s1_reset_n <= reset_n;
  gen_code_value_pio_0_s1_chipselect <= internal_nios2_clock_6_out_granted_gen_code_value_pio_0_s1;
  --gen_code_value_pio_0_s1_firsttransfer first transaction, which is an e_assign
  gen_code_value_pio_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(gen_code_value_pio_0_s1_begins_xfer) = '1'), gen_code_value_pio_0_s1_unreg_firsttransfer, gen_code_value_pio_0_s1_reg_firsttransfer);
  --gen_code_value_pio_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  gen_code_value_pio_0_s1_unreg_firsttransfer <= NOT ((gen_code_value_pio_0_s1_slavearbiterlockenable AND gen_code_value_pio_0_s1_any_continuerequest));
  --gen_code_value_pio_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_value_pio_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gen_code_value_pio_0_s1_begins_xfer) = '1' then 
        gen_code_value_pio_0_s1_reg_firsttransfer <= gen_code_value_pio_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gen_code_value_pio_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gen_code_value_pio_0_s1_beginbursttransfer_internal <= gen_code_value_pio_0_s1_begins_xfer;
  --~gen_code_value_pio_0_s1_write_n assignment, which is an e_mux
  gen_code_value_pio_0_s1_write_n <= NOT ((internal_nios2_clock_6_out_granted_gen_code_value_pio_0_s1 AND nios2_clock_6_out_write));
  --gen_code_value_pio_0_s1_address mux, which is an e_mux
  gen_code_value_pio_0_s1_address <= nios2_clock_6_out_nativeaddress;
  --d1_gen_code_value_pio_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gen_code_value_pio_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gen_code_value_pio_0_s1_end_xfer <= gen_code_value_pio_0_s1_end_xfer;
    end if;

  end process;

  --gen_code_value_pio_0_s1_waits_for_read in a cycle, which is an e_mux
  gen_code_value_pio_0_s1_waits_for_read <= gen_code_value_pio_0_s1_in_a_read_cycle AND gen_code_value_pio_0_s1_begins_xfer;
  --gen_code_value_pio_0_s1_in_a_read_cycle assignment, which is an e_assign
  gen_code_value_pio_0_s1_in_a_read_cycle <= internal_nios2_clock_6_out_granted_gen_code_value_pio_0_s1 AND nios2_clock_6_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gen_code_value_pio_0_s1_in_a_read_cycle;
  --gen_code_value_pio_0_s1_waits_for_write in a cycle, which is an e_mux
  gen_code_value_pio_0_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_value_pio_0_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --gen_code_value_pio_0_s1_in_a_write_cycle assignment, which is an e_assign
  gen_code_value_pio_0_s1_in_a_write_cycle <= internal_nios2_clock_6_out_granted_gen_code_value_pio_0_s1 AND nios2_clock_6_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gen_code_value_pio_0_s1_in_a_write_cycle;
  wait_for_gen_code_value_pio_0_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_6_out_granted_gen_code_value_pio_0_s1 <= internal_nios2_clock_6_out_granted_gen_code_value_pio_0_s1;
  --vhdl renameroo for output signals
  nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 <= internal_nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1;
  --vhdl renameroo for output signals
  nios2_clock_6_out_requests_gen_code_value_pio_0_s1 <= internal_nios2_clock_6_out_requests_gen_code_value_pio_0_s1;
--synthesis translate_off
    --gen_code_value_pio_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gen_code_value_pio_1_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal gen_code_value_pio_1_s1_readdata : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal nios2_clock_7_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_7_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_7_out_read : IN STD_LOGIC;
                 signal nios2_clock_7_out_write : IN STD_LOGIC;
                 signal nios2_clock_7_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_gen_code_value_pio_1_s1_end_xfer : OUT STD_LOGIC;
                 signal gen_code_value_pio_1_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gen_code_value_pio_1_s1_chipselect : OUT STD_LOGIC;
                 signal gen_code_value_pio_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal gen_code_value_pio_1_s1_reset_n : OUT STD_LOGIC;
                 signal gen_code_value_pio_1_s1_write_n : OUT STD_LOGIC;
                 signal gen_code_value_pio_1_s1_writedata : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal nios2_clock_7_out_granted_gen_code_value_pio_1_s1 : OUT STD_LOGIC;
                 signal nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 : OUT STD_LOGIC;
                 signal nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1 : OUT STD_LOGIC;
                 signal nios2_clock_7_out_requests_gen_code_value_pio_1_s1 : OUT STD_LOGIC
              );
end entity gen_code_value_pio_1_s1_arbitrator;


architecture europa of gen_code_value_pio_1_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_allgrants :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_any_continuerequest :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_arb_counter_enable :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_arb_share_counter :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_arb_share_set_values :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_begins_xfer :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_end_xfer :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_firsttransfer :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_grant_vector :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_in_a_read_cycle :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_in_a_write_cycle :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_master_qreq_vector :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_non_bursting_master_requests :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_reg_firsttransfer :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_slavearbiterlockenable :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_unreg_firsttransfer :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_waits_for_read :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_7_out_granted_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal internal_nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal internal_nios2_clock_7_out_requests_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal nios2_clock_7_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_7_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_7_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_7_out_saved_grant_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal wait_for_gen_code_value_pio_1_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gen_code_value_pio_1_s1_end_xfer;
    end if;

  end process;

  gen_code_value_pio_1_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1);
  --assign gen_code_value_pio_1_s1_readdata_from_sa = gen_code_value_pio_1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gen_code_value_pio_1_s1_readdata_from_sa <= gen_code_value_pio_1_s1_readdata;
  internal_nios2_clock_7_out_requests_gen_code_value_pio_1_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_7_out_read OR nios2_clock_7_out_write)))))));
  --gen_code_value_pio_1_s1_arb_share_counter set values, which is an e_mux
  gen_code_value_pio_1_s1_arb_share_set_values <= std_logic'('1');
  --gen_code_value_pio_1_s1_non_bursting_master_requests mux, which is an e_mux
  gen_code_value_pio_1_s1_non_bursting_master_requests <= internal_nios2_clock_7_out_requests_gen_code_value_pio_1_s1;
  --gen_code_value_pio_1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  gen_code_value_pio_1_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --gen_code_value_pio_1_s1_arb_share_counter_next_value assignment, which is an e_assign
  gen_code_value_pio_1_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gen_code_value_pio_1_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_value_pio_1_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gen_code_value_pio_1_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_value_pio_1_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gen_code_value_pio_1_s1_allgrants all slave grants, which is an e_mux
  gen_code_value_pio_1_s1_allgrants <= gen_code_value_pio_1_s1_grant_vector;
  --gen_code_value_pio_1_s1_end_xfer assignment, which is an e_assign
  gen_code_value_pio_1_s1_end_xfer <= NOT ((gen_code_value_pio_1_s1_waits_for_read OR gen_code_value_pio_1_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_gen_code_value_pio_1_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gen_code_value_pio_1_s1 <= gen_code_value_pio_1_s1_end_xfer AND (((NOT gen_code_value_pio_1_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gen_code_value_pio_1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  gen_code_value_pio_1_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gen_code_value_pio_1_s1 AND gen_code_value_pio_1_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_gen_code_value_pio_1_s1 AND NOT gen_code_value_pio_1_s1_non_bursting_master_requests));
  --gen_code_value_pio_1_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_value_pio_1_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gen_code_value_pio_1_s1_arb_counter_enable) = '1' then 
        gen_code_value_pio_1_s1_arb_share_counter <= gen_code_value_pio_1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gen_code_value_pio_1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_value_pio_1_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gen_code_value_pio_1_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_gen_code_value_pio_1_s1)) OR ((end_xfer_arb_share_counter_term_gen_code_value_pio_1_s1 AND NOT gen_code_value_pio_1_s1_non_bursting_master_requests)))) = '1' then 
        gen_code_value_pio_1_s1_slavearbiterlockenable <= gen_code_value_pio_1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_7/out gen_code_value_pio_1/s1 arbiterlock, which is an e_assign
  nios2_clock_7_out_arbiterlock <= gen_code_value_pio_1_s1_slavearbiterlockenable AND nios2_clock_7_out_continuerequest;
  --gen_code_value_pio_1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gen_code_value_pio_1_s1_slavearbiterlockenable2 <= gen_code_value_pio_1_s1_arb_share_counter_next_value;
  --nios2_clock_7/out gen_code_value_pio_1/s1 arbiterlock2, which is an e_assign
  nios2_clock_7_out_arbiterlock2 <= gen_code_value_pio_1_s1_slavearbiterlockenable2 AND nios2_clock_7_out_continuerequest;
  --gen_code_value_pio_1_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  gen_code_value_pio_1_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_7_out_continuerequest continued request, which is an e_assign
  nios2_clock_7_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 <= internal_nios2_clock_7_out_requests_gen_code_value_pio_1_s1;
  --gen_code_value_pio_1_s1_writedata mux, which is an e_mux
  gen_code_value_pio_1_s1_writedata <= nios2_clock_7_out_writedata (23 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_clock_7_out_granted_gen_code_value_pio_1_s1 <= internal_nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1;
  --nios2_clock_7/out saved-grant gen_code_value_pio_1/s1, which is an e_assign
  nios2_clock_7_out_saved_grant_gen_code_value_pio_1_s1 <= internal_nios2_clock_7_out_requests_gen_code_value_pio_1_s1;
  --allow new arb cycle for gen_code_value_pio_1/s1, which is an e_assign
  gen_code_value_pio_1_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gen_code_value_pio_1_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gen_code_value_pio_1_s1_master_qreq_vector <= std_logic'('1');
  --gen_code_value_pio_1_s1_reset_n assignment, which is an e_assign
  gen_code_value_pio_1_s1_reset_n <= reset_n;
  gen_code_value_pio_1_s1_chipselect <= internal_nios2_clock_7_out_granted_gen_code_value_pio_1_s1;
  --gen_code_value_pio_1_s1_firsttransfer first transaction, which is an e_assign
  gen_code_value_pio_1_s1_firsttransfer <= A_WE_StdLogic((std_logic'(gen_code_value_pio_1_s1_begins_xfer) = '1'), gen_code_value_pio_1_s1_unreg_firsttransfer, gen_code_value_pio_1_s1_reg_firsttransfer);
  --gen_code_value_pio_1_s1_unreg_firsttransfer first transaction, which is an e_assign
  gen_code_value_pio_1_s1_unreg_firsttransfer <= NOT ((gen_code_value_pio_1_s1_slavearbiterlockenable AND gen_code_value_pio_1_s1_any_continuerequest));
  --gen_code_value_pio_1_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gen_code_value_pio_1_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gen_code_value_pio_1_s1_begins_xfer) = '1' then 
        gen_code_value_pio_1_s1_reg_firsttransfer <= gen_code_value_pio_1_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gen_code_value_pio_1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gen_code_value_pio_1_s1_beginbursttransfer_internal <= gen_code_value_pio_1_s1_begins_xfer;
  --~gen_code_value_pio_1_s1_write_n assignment, which is an e_mux
  gen_code_value_pio_1_s1_write_n <= NOT ((internal_nios2_clock_7_out_granted_gen_code_value_pio_1_s1 AND nios2_clock_7_out_write));
  --gen_code_value_pio_1_s1_address mux, which is an e_mux
  gen_code_value_pio_1_s1_address <= nios2_clock_7_out_nativeaddress;
  --d1_gen_code_value_pio_1_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gen_code_value_pio_1_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gen_code_value_pio_1_s1_end_xfer <= gen_code_value_pio_1_s1_end_xfer;
    end if;

  end process;

  --gen_code_value_pio_1_s1_waits_for_read in a cycle, which is an e_mux
  gen_code_value_pio_1_s1_waits_for_read <= gen_code_value_pio_1_s1_in_a_read_cycle AND gen_code_value_pio_1_s1_begins_xfer;
  --gen_code_value_pio_1_s1_in_a_read_cycle assignment, which is an e_assign
  gen_code_value_pio_1_s1_in_a_read_cycle <= internal_nios2_clock_7_out_granted_gen_code_value_pio_1_s1 AND nios2_clock_7_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gen_code_value_pio_1_s1_in_a_read_cycle;
  --gen_code_value_pio_1_s1_waits_for_write in a cycle, which is an e_mux
  gen_code_value_pio_1_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gen_code_value_pio_1_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --gen_code_value_pio_1_s1_in_a_write_cycle assignment, which is an e_assign
  gen_code_value_pio_1_s1_in_a_write_cycle <= internal_nios2_clock_7_out_granted_gen_code_value_pio_1_s1 AND nios2_clock_7_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gen_code_value_pio_1_s1_in_a_write_cycle;
  wait_for_gen_code_value_pio_1_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_7_out_granted_gen_code_value_pio_1_s1 <= internal_nios2_clock_7_out_granted_gen_code_value_pio_1_s1;
  --vhdl renameroo for output signals
  nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 <= internal_nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1;
  --vhdl renameroo for output signals
  nios2_clock_7_out_requests_gen_code_value_pio_1_s1 <= internal_nios2_clock_7_out_requests_gen_code_value_pio_1_s1;
--synthesis translate_off
    --gen_code_value_pio_1/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_0_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_0_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal nios2_clock_2_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_2_out_nativeaddress : IN STD_LOGIC;
                 signal nios2_clock_2_out_read : IN STD_LOGIC;
                 signal nios2_clock_2_out_write : IN STD_LOGIC;
                 signal nios2_clock_2_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                 signal nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                 signal nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                 signal nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC
              );
end entity jtag_uart_0_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_0_avalon_jtag_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal internal_nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal internal_nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_share_counter :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal nios2_clock_2_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_2_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_2_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_2_out_saved_grant_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal wait_for_jtag_uart_0_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_0_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_0_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave);
  --assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_readdata_from_sa <= jtag_uart_0_avalon_jtag_slave_readdata;
  internal_nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_2_out_read OR nios2_clock_2_out_write)))))));
  --assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_0_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_0_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_0_avalon_jtag_slave_waitrequest;
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_arb_share_set_values <= std_logic'('1');
  --jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests <= internal_nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave;
  --jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(jtag_uart_0_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_0_avalon_jtag_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(jtag_uart_0_avalon_jtag_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_0_avalon_jtag_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --jtag_uart_0_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_allgrants <= jtag_uart_0_avalon_jtag_slave_grant_vector;
  --jtag_uart_0_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_0_avalon_jtag_slave_waits_for_read OR jtag_uart_0_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave <= jtag_uart_0_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave AND jtag_uart_0_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave AND NOT jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_0_avalon_jtag_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_0_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_0_avalon_jtag_slave_arb_share_counter <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_0_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave AND NOT jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_2/out jtag_uart_0/avalon_jtag_slave arbiterlock, which is an e_assign
  nios2_clock_2_out_arbiterlock <= jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable AND nios2_clock_2_out_continuerequest;
  --jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
  --nios2_clock_2/out jtag_uart_0/avalon_jtag_slave arbiterlock2, which is an e_assign
  nios2_clock_2_out_arbiterlock2 <= jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 AND nios2_clock_2_out_continuerequest;
  --jtag_uart_0_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --nios2_clock_2_out_continuerequest continued request, which is an e_assign
  nios2_clock_2_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave <= internal_nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave;
  --jtag_uart_0_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_writedata <= nios2_clock_2_out_writedata;
  --master is always granted when requested
  internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave <= internal_nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave;
  --nios2_clock_2/out saved-grant jtag_uart_0/avalon_jtag_slave, which is an e_assign
  nios2_clock_2_out_saved_grant_jtag_uart_0_avalon_jtag_slave <= internal_nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart_0/avalon_jtag_slave, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_0_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_0_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_0_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_0_avalon_jtag_slave_chipselect <= internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave;
  --jtag_uart_0_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_0_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_0_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_0_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_0_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_0_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_0_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_0_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_read_n <= NOT ((internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave AND nios2_clock_2_out_read));
  --~jtag_uart_0_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_write_n <= NOT ((internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave AND nios2_clock_2_out_write));
  --jtag_uart_0_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_address <= nios2_clock_2_out_nativeaddress;
  --d1_jtag_uart_0_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= jtag_uart_0_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_0_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_waits_for_read <= jtag_uart_0_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_0_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_in_a_read_cycle <= internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave AND nios2_clock_2_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_0_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_waits_for_write <= jtag_uart_0_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_0_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_in_a_write_cycle <= internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave AND nios2_clock_2_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_0_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_irq_from_sa <= jtag_uart_0_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave <= internal_nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave;
  --vhdl renameroo for output signals
  nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave <= internal_nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave;
  --vhdl renameroo for output signals
  nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave <= internal_nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave;
--synthesis translate_off
    --jtag_uart_0/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity latch_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal latch_pio_s1_readdata : IN STD_LOGIC;
                 signal nios2_clock_18_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_18_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_18_out_read : IN STD_LOGIC;
                 signal nios2_clock_18_out_write : IN STD_LOGIC;
                 signal nios2_clock_18_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_latch_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal latch_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal latch_pio_s1_chipselect : OUT STD_LOGIC;
                 signal latch_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal latch_pio_s1_reset_n : OUT STD_LOGIC;
                 signal latch_pio_s1_write_n : OUT STD_LOGIC;
                 signal latch_pio_s1_writedata : OUT STD_LOGIC;
                 signal nios2_clock_18_out_granted_latch_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_18_out_qualified_request_latch_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_18_out_read_data_valid_latch_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_18_out_requests_latch_pio_s1 : OUT STD_LOGIC
              );
end entity latch_pio_s1_arbitrator;


architecture europa of latch_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_latch_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_18_out_granted_latch_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_18_out_qualified_request_latch_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_18_out_requests_latch_pio_s1 :  STD_LOGIC;
                signal latch_pio_s1_allgrants :  STD_LOGIC;
                signal latch_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal latch_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal latch_pio_s1_any_continuerequest :  STD_LOGIC;
                signal latch_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal latch_pio_s1_arb_share_counter :  STD_LOGIC;
                signal latch_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal latch_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal latch_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal latch_pio_s1_begins_xfer :  STD_LOGIC;
                signal latch_pio_s1_end_xfer :  STD_LOGIC;
                signal latch_pio_s1_firsttransfer :  STD_LOGIC;
                signal latch_pio_s1_grant_vector :  STD_LOGIC;
                signal latch_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal latch_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal latch_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal latch_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal latch_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal latch_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal latch_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal latch_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal latch_pio_s1_waits_for_read :  STD_LOGIC;
                signal latch_pio_s1_waits_for_write :  STD_LOGIC;
                signal nios2_clock_18_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_18_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_18_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_18_out_saved_grant_latch_pio_s1 :  STD_LOGIC;
                signal wait_for_latch_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT latch_pio_s1_end_xfer;
    end if;

  end process;

  latch_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_18_out_qualified_request_latch_pio_s1);
  --assign latch_pio_s1_readdata_from_sa = latch_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  latch_pio_s1_readdata_from_sa <= latch_pio_s1_readdata;
  internal_nios2_clock_18_out_requests_latch_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_18_out_read OR nios2_clock_18_out_write)))))));
  --latch_pio_s1_arb_share_counter set values, which is an e_mux
  latch_pio_s1_arb_share_set_values <= std_logic'('1');
  --latch_pio_s1_non_bursting_master_requests mux, which is an e_mux
  latch_pio_s1_non_bursting_master_requests <= internal_nios2_clock_18_out_requests_latch_pio_s1;
  --latch_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  latch_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --latch_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  latch_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(latch_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latch_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(latch_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latch_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --latch_pio_s1_allgrants all slave grants, which is an e_mux
  latch_pio_s1_allgrants <= latch_pio_s1_grant_vector;
  --latch_pio_s1_end_xfer assignment, which is an e_assign
  latch_pio_s1_end_xfer <= NOT ((latch_pio_s1_waits_for_read OR latch_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_latch_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_latch_pio_s1 <= latch_pio_s1_end_xfer AND (((NOT latch_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --latch_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  latch_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_latch_pio_s1 AND latch_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_latch_pio_s1 AND NOT latch_pio_s1_non_bursting_master_requests));
  --latch_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      latch_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(latch_pio_s1_arb_counter_enable) = '1' then 
        latch_pio_s1_arb_share_counter <= latch_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --latch_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      latch_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((latch_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_latch_pio_s1)) OR ((end_xfer_arb_share_counter_term_latch_pio_s1 AND NOT latch_pio_s1_non_bursting_master_requests)))) = '1' then 
        latch_pio_s1_slavearbiterlockenable <= latch_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_18/out latch_pio/s1 arbiterlock, which is an e_assign
  nios2_clock_18_out_arbiterlock <= latch_pio_s1_slavearbiterlockenable AND nios2_clock_18_out_continuerequest;
  --latch_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  latch_pio_s1_slavearbiterlockenable2 <= latch_pio_s1_arb_share_counter_next_value;
  --nios2_clock_18/out latch_pio/s1 arbiterlock2, which is an e_assign
  nios2_clock_18_out_arbiterlock2 <= latch_pio_s1_slavearbiterlockenable2 AND nios2_clock_18_out_continuerequest;
  --latch_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  latch_pio_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_18_out_continuerequest continued request, which is an e_assign
  nios2_clock_18_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_18_out_qualified_request_latch_pio_s1 <= internal_nios2_clock_18_out_requests_latch_pio_s1;
  --latch_pio_s1_writedata mux, which is an e_mux
  latch_pio_s1_writedata <= nios2_clock_18_out_writedata(0);
  --master is always granted when requested
  internal_nios2_clock_18_out_granted_latch_pio_s1 <= internal_nios2_clock_18_out_qualified_request_latch_pio_s1;
  --nios2_clock_18/out saved-grant latch_pio/s1, which is an e_assign
  nios2_clock_18_out_saved_grant_latch_pio_s1 <= internal_nios2_clock_18_out_requests_latch_pio_s1;
  --allow new arb cycle for latch_pio/s1, which is an e_assign
  latch_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  latch_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  latch_pio_s1_master_qreq_vector <= std_logic'('1');
  --latch_pio_s1_reset_n assignment, which is an e_assign
  latch_pio_s1_reset_n <= reset_n;
  latch_pio_s1_chipselect <= internal_nios2_clock_18_out_granted_latch_pio_s1;
  --latch_pio_s1_firsttransfer first transaction, which is an e_assign
  latch_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(latch_pio_s1_begins_xfer) = '1'), latch_pio_s1_unreg_firsttransfer, latch_pio_s1_reg_firsttransfer);
  --latch_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  latch_pio_s1_unreg_firsttransfer <= NOT ((latch_pio_s1_slavearbiterlockenable AND latch_pio_s1_any_continuerequest));
  --latch_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      latch_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(latch_pio_s1_begins_xfer) = '1' then 
        latch_pio_s1_reg_firsttransfer <= latch_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --latch_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  latch_pio_s1_beginbursttransfer_internal <= latch_pio_s1_begins_xfer;
  --~latch_pio_s1_write_n assignment, which is an e_mux
  latch_pio_s1_write_n <= NOT ((internal_nios2_clock_18_out_granted_latch_pio_s1 AND nios2_clock_18_out_write));
  --latch_pio_s1_address mux, which is an e_mux
  latch_pio_s1_address <= nios2_clock_18_out_nativeaddress;
  --d1_latch_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_latch_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_latch_pio_s1_end_xfer <= latch_pio_s1_end_xfer;
    end if;

  end process;

  --latch_pio_s1_waits_for_read in a cycle, which is an e_mux
  latch_pio_s1_waits_for_read <= latch_pio_s1_in_a_read_cycle AND latch_pio_s1_begins_xfer;
  --latch_pio_s1_in_a_read_cycle assignment, which is an e_assign
  latch_pio_s1_in_a_read_cycle <= internal_nios2_clock_18_out_granted_latch_pio_s1 AND nios2_clock_18_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= latch_pio_s1_in_a_read_cycle;
  --latch_pio_s1_waits_for_write in a cycle, which is an e_mux
  latch_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latch_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --latch_pio_s1_in_a_write_cycle assignment, which is an e_assign
  latch_pio_s1_in_a_write_cycle <= internal_nios2_clock_18_out_granted_latch_pio_s1 AND nios2_clock_18_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= latch_pio_s1_in_a_write_cycle;
  wait_for_latch_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_18_out_granted_latch_pio_s1 <= internal_nios2_clock_18_out_granted_latch_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_18_out_qualified_request_latch_pio_s1 <= internal_nios2_clock_18_out_qualified_request_latch_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_18_out_requests_latch_pio_s1 <= internal_nios2_clock_18_out_requests_latch_pio_s1;
--synthesis translate_off
    --latch_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity led_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_12_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_12_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_12_out_read : IN STD_LOGIC;
                 signal nios2_clock_12_out_write : IN STD_LOGIC;
                 signal nios2_clock_12_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal led_pio_s1_chipselect : OUT STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal led_pio_s1_reset_n : OUT STD_LOGIC;
                 signal led_pio_s1_write_n : OUT STD_LOGIC;
                 signal led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_12_out_granted_led_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_12_out_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_12_out_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_12_out_requests_led_pio_s1 : OUT STD_LOGIC
              );
end entity led_pio_s1_arbitrator;


architecture europa of led_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_led_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_12_out_granted_led_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_12_out_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_12_out_requests_led_pio_s1 :  STD_LOGIC;
                signal led_pio_s1_allgrants :  STD_LOGIC;
                signal led_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal led_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal led_pio_s1_any_continuerequest :  STD_LOGIC;
                signal led_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal led_pio_s1_arb_share_counter :  STD_LOGIC;
                signal led_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal led_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal led_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal led_pio_s1_begins_xfer :  STD_LOGIC;
                signal led_pio_s1_end_xfer :  STD_LOGIC;
                signal led_pio_s1_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_grant_vector :  STD_LOGIC;
                signal led_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal led_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal led_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal led_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal led_pio_s1_pretend_byte_enable :  STD_LOGIC;
                signal led_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal led_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_waits_for_read :  STD_LOGIC;
                signal led_pio_s1_waits_for_write :  STD_LOGIC;
                signal nios2_clock_12_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_12_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_12_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_12_out_saved_grant_led_pio_s1 :  STD_LOGIC;
                signal wait_for_led_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT led_pio_s1_end_xfer;
    end if;

  end process;

  led_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_12_out_qualified_request_led_pio_s1);
  --assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  led_pio_s1_readdata_from_sa <= led_pio_s1_readdata;
  internal_nios2_clock_12_out_requests_led_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_12_out_read OR nios2_clock_12_out_write)))))));
  --led_pio_s1_arb_share_counter set values, which is an e_mux
  led_pio_s1_arb_share_set_values <= std_logic'('1');
  --led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  led_pio_s1_non_bursting_master_requests <= internal_nios2_clock_12_out_requests_led_pio_s1;
  --led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  led_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  led_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(led_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(led_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --led_pio_s1_allgrants all slave grants, which is an e_mux
  led_pio_s1_allgrants <= led_pio_s1_grant_vector;
  --led_pio_s1_end_xfer assignment, which is an e_assign
  led_pio_s1_end_xfer <= NOT ((led_pio_s1_waits_for_read OR led_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_led_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_led_pio_s1 <= led_pio_s1_end_xfer AND (((NOT led_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  led_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_led_pio_s1 AND led_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests));
  --led_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_arb_counter_enable) = '1' then 
        led_pio_s1_arb_share_counter <= led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((led_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_led_pio_s1)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests)))) = '1' then 
        led_pio_s1_slavearbiterlockenable <= led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_12/out led_pio/s1 arbiterlock, which is an e_assign
  nios2_clock_12_out_arbiterlock <= led_pio_s1_slavearbiterlockenable AND nios2_clock_12_out_continuerequest;
  --led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  led_pio_s1_slavearbiterlockenable2 <= led_pio_s1_arb_share_counter_next_value;
  --nios2_clock_12/out led_pio/s1 arbiterlock2, which is an e_assign
  nios2_clock_12_out_arbiterlock2 <= led_pio_s1_slavearbiterlockenable2 AND nios2_clock_12_out_continuerequest;
  --led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  led_pio_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_12_out_continuerequest continued request, which is an e_assign
  nios2_clock_12_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_12_out_qualified_request_led_pio_s1 <= internal_nios2_clock_12_out_requests_led_pio_s1;
  --led_pio_s1_writedata mux, which is an e_mux
  led_pio_s1_writedata <= nios2_clock_12_out_writedata;
  --master is always granted when requested
  internal_nios2_clock_12_out_granted_led_pio_s1 <= internal_nios2_clock_12_out_qualified_request_led_pio_s1;
  --nios2_clock_12/out saved-grant led_pio/s1, which is an e_assign
  nios2_clock_12_out_saved_grant_led_pio_s1 <= internal_nios2_clock_12_out_requests_led_pio_s1;
  --allow new arb cycle for led_pio/s1, which is an e_assign
  led_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  led_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  led_pio_s1_master_qreq_vector <= std_logic'('1');
  --led_pio_s1_reset_n assignment, which is an e_assign
  led_pio_s1_reset_n <= reset_n;
  led_pio_s1_chipselect <= internal_nios2_clock_12_out_granted_led_pio_s1;
  --led_pio_s1_firsttransfer first transaction, which is an e_assign
  led_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(led_pio_s1_begins_xfer) = '1'), led_pio_s1_unreg_firsttransfer, led_pio_s1_reg_firsttransfer);
  --led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  led_pio_s1_unreg_firsttransfer <= NOT ((led_pio_s1_slavearbiterlockenable AND led_pio_s1_any_continuerequest));
  --led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_begins_xfer) = '1' then 
        led_pio_s1_reg_firsttransfer <= led_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  led_pio_s1_beginbursttransfer_internal <= led_pio_s1_begins_xfer;
  --~led_pio_s1_write_n assignment, which is an e_mux
  led_pio_s1_write_n <= NOT ((((internal_nios2_clock_12_out_granted_led_pio_s1 AND nios2_clock_12_out_write)) AND led_pio_s1_pretend_byte_enable));
  --led_pio_s1_address mux, which is an e_mux
  led_pio_s1_address <= nios2_clock_12_out_nativeaddress;
  --d1_led_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_led_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_led_pio_s1_end_xfer <= led_pio_s1_end_xfer;
    end if;

  end process;

  --led_pio_s1_waits_for_read in a cycle, which is an e_mux
  led_pio_s1_waits_for_read <= led_pio_s1_in_a_read_cycle AND led_pio_s1_begins_xfer;
  --led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  led_pio_s1_in_a_read_cycle <= internal_nios2_clock_12_out_granted_led_pio_s1 AND nios2_clock_12_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= led_pio_s1_in_a_read_cycle;
  --led_pio_s1_waits_for_write in a cycle, which is an e_mux
  led_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  led_pio_s1_in_a_write_cycle <= internal_nios2_clock_12_out_granted_led_pio_s1 AND nios2_clock_12_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= led_pio_s1_in_a_write_cycle;
  wait_for_led_pio_s1_counter <= std_logic'('0');
  --led_pio_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  led_pio_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_nios2_clock_12_out_granted_led_pio_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(std_logic'('1')))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  nios2_clock_12_out_granted_led_pio_s1 <= internal_nios2_clock_12_out_granted_led_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_12_out_qualified_request_led_pio_s1 <= internal_nios2_clock_12_out_qualified_request_led_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_12_out_requests_led_pio_s1 <= internal_nios2_clock_12_out_requests_led_pio_s1;
--synthesis translate_off
    --led_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity mode_select_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal mode_select_s1_readdata : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_out_read : IN STD_LOGIC;
                 signal nios2_clock_10_out_write : IN STD_LOGIC;
                 signal nios2_clock_10_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_mode_select_s1_end_xfer : OUT STD_LOGIC;
                 signal mode_select_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mode_select_s1_chipselect : OUT STD_LOGIC;
                 signal mode_select_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mode_select_s1_reset_n : OUT STD_LOGIC;
                 signal mode_select_s1_write_n : OUT STD_LOGIC;
                 signal mode_select_s1_writedata : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_out_granted_mode_select_s1 : OUT STD_LOGIC;
                 signal nios2_clock_10_out_qualified_request_mode_select_s1 : OUT STD_LOGIC;
                 signal nios2_clock_10_out_read_data_valid_mode_select_s1 : OUT STD_LOGIC;
                 signal nios2_clock_10_out_requests_mode_select_s1 : OUT STD_LOGIC
              );
end entity mode_select_s1_arbitrator;


architecture europa of mode_select_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_mode_select_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_10_out_granted_mode_select_s1 :  STD_LOGIC;
                signal internal_nios2_clock_10_out_qualified_request_mode_select_s1 :  STD_LOGIC;
                signal internal_nios2_clock_10_out_requests_mode_select_s1 :  STD_LOGIC;
                signal mode_select_s1_allgrants :  STD_LOGIC;
                signal mode_select_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal mode_select_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal mode_select_s1_any_continuerequest :  STD_LOGIC;
                signal mode_select_s1_arb_counter_enable :  STD_LOGIC;
                signal mode_select_s1_arb_share_counter :  STD_LOGIC;
                signal mode_select_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal mode_select_s1_arb_share_set_values :  STD_LOGIC;
                signal mode_select_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal mode_select_s1_begins_xfer :  STD_LOGIC;
                signal mode_select_s1_end_xfer :  STD_LOGIC;
                signal mode_select_s1_firsttransfer :  STD_LOGIC;
                signal mode_select_s1_grant_vector :  STD_LOGIC;
                signal mode_select_s1_in_a_read_cycle :  STD_LOGIC;
                signal mode_select_s1_in_a_write_cycle :  STD_LOGIC;
                signal mode_select_s1_master_qreq_vector :  STD_LOGIC;
                signal mode_select_s1_non_bursting_master_requests :  STD_LOGIC;
                signal mode_select_s1_reg_firsttransfer :  STD_LOGIC;
                signal mode_select_s1_slavearbiterlockenable :  STD_LOGIC;
                signal mode_select_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal mode_select_s1_unreg_firsttransfer :  STD_LOGIC;
                signal mode_select_s1_waits_for_read :  STD_LOGIC;
                signal mode_select_s1_waits_for_write :  STD_LOGIC;
                signal nios2_clock_10_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_10_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_10_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_10_out_saved_grant_mode_select_s1 :  STD_LOGIC;
                signal wait_for_mode_select_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT mode_select_s1_end_xfer;
    end if;

  end process;

  mode_select_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_10_out_qualified_request_mode_select_s1);
  --assign mode_select_s1_readdata_from_sa = mode_select_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  mode_select_s1_readdata_from_sa <= mode_select_s1_readdata;
  internal_nios2_clock_10_out_requests_mode_select_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_10_out_read OR nios2_clock_10_out_write)))))));
  --mode_select_s1_arb_share_counter set values, which is an e_mux
  mode_select_s1_arb_share_set_values <= std_logic'('1');
  --mode_select_s1_non_bursting_master_requests mux, which is an e_mux
  mode_select_s1_non_bursting_master_requests <= internal_nios2_clock_10_out_requests_mode_select_s1;
  --mode_select_s1_any_bursting_master_saved_grant mux, which is an e_mux
  mode_select_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --mode_select_s1_arb_share_counter_next_value assignment, which is an e_assign
  mode_select_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(mode_select_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mode_select_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(mode_select_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mode_select_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --mode_select_s1_allgrants all slave grants, which is an e_mux
  mode_select_s1_allgrants <= mode_select_s1_grant_vector;
  --mode_select_s1_end_xfer assignment, which is an e_assign
  mode_select_s1_end_xfer <= NOT ((mode_select_s1_waits_for_read OR mode_select_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_mode_select_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_mode_select_s1 <= mode_select_s1_end_xfer AND (((NOT mode_select_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --mode_select_s1_arb_share_counter arbitration counter enable, which is an e_assign
  mode_select_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_mode_select_s1 AND mode_select_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_mode_select_s1 AND NOT mode_select_s1_non_bursting_master_requests));
  --mode_select_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      mode_select_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(mode_select_s1_arb_counter_enable) = '1' then 
        mode_select_s1_arb_share_counter <= mode_select_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --mode_select_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      mode_select_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((mode_select_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_mode_select_s1)) OR ((end_xfer_arb_share_counter_term_mode_select_s1 AND NOT mode_select_s1_non_bursting_master_requests)))) = '1' then 
        mode_select_s1_slavearbiterlockenable <= mode_select_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_10/out mode_select/s1 arbiterlock, which is an e_assign
  nios2_clock_10_out_arbiterlock <= mode_select_s1_slavearbiterlockenable AND nios2_clock_10_out_continuerequest;
  --mode_select_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  mode_select_s1_slavearbiterlockenable2 <= mode_select_s1_arb_share_counter_next_value;
  --nios2_clock_10/out mode_select/s1 arbiterlock2, which is an e_assign
  nios2_clock_10_out_arbiterlock2 <= mode_select_s1_slavearbiterlockenable2 AND nios2_clock_10_out_continuerequest;
  --mode_select_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  mode_select_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_10_out_continuerequest continued request, which is an e_assign
  nios2_clock_10_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_10_out_qualified_request_mode_select_s1 <= internal_nios2_clock_10_out_requests_mode_select_s1;
  --mode_select_s1_writedata mux, which is an e_mux
  mode_select_s1_writedata <= nios2_clock_10_out_writedata (1 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_clock_10_out_granted_mode_select_s1 <= internal_nios2_clock_10_out_qualified_request_mode_select_s1;
  --nios2_clock_10/out saved-grant mode_select/s1, which is an e_assign
  nios2_clock_10_out_saved_grant_mode_select_s1 <= internal_nios2_clock_10_out_requests_mode_select_s1;
  --allow new arb cycle for mode_select/s1, which is an e_assign
  mode_select_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  mode_select_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  mode_select_s1_master_qreq_vector <= std_logic'('1');
  --mode_select_s1_reset_n assignment, which is an e_assign
  mode_select_s1_reset_n <= reset_n;
  mode_select_s1_chipselect <= internal_nios2_clock_10_out_granted_mode_select_s1;
  --mode_select_s1_firsttransfer first transaction, which is an e_assign
  mode_select_s1_firsttransfer <= A_WE_StdLogic((std_logic'(mode_select_s1_begins_xfer) = '1'), mode_select_s1_unreg_firsttransfer, mode_select_s1_reg_firsttransfer);
  --mode_select_s1_unreg_firsttransfer first transaction, which is an e_assign
  mode_select_s1_unreg_firsttransfer <= NOT ((mode_select_s1_slavearbiterlockenable AND mode_select_s1_any_continuerequest));
  --mode_select_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      mode_select_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(mode_select_s1_begins_xfer) = '1' then 
        mode_select_s1_reg_firsttransfer <= mode_select_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --mode_select_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  mode_select_s1_beginbursttransfer_internal <= mode_select_s1_begins_xfer;
  --~mode_select_s1_write_n assignment, which is an e_mux
  mode_select_s1_write_n <= NOT ((internal_nios2_clock_10_out_granted_mode_select_s1 AND nios2_clock_10_out_write));
  --mode_select_s1_address mux, which is an e_mux
  mode_select_s1_address <= nios2_clock_10_out_nativeaddress;
  --d1_mode_select_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_mode_select_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_mode_select_s1_end_xfer <= mode_select_s1_end_xfer;
    end if;

  end process;

  --mode_select_s1_waits_for_read in a cycle, which is an e_mux
  mode_select_s1_waits_for_read <= mode_select_s1_in_a_read_cycle AND mode_select_s1_begins_xfer;
  --mode_select_s1_in_a_read_cycle assignment, which is an e_assign
  mode_select_s1_in_a_read_cycle <= internal_nios2_clock_10_out_granted_mode_select_s1 AND nios2_clock_10_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= mode_select_s1_in_a_read_cycle;
  --mode_select_s1_waits_for_write in a cycle, which is an e_mux
  mode_select_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mode_select_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --mode_select_s1_in_a_write_cycle assignment, which is an e_assign
  mode_select_s1_in_a_write_cycle <= internal_nios2_clock_10_out_granted_mode_select_s1 AND nios2_clock_10_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= mode_select_s1_in_a_write_cycle;
  wait_for_mode_select_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_10_out_granted_mode_select_s1 <= internal_nios2_clock_10_out_granted_mode_select_s1;
  --vhdl renameroo for output signals
  nios2_clock_10_out_qualified_request_mode_select_s1 <= internal_nios2_clock_10_out_qualified_request_mode_select_s1;
  --vhdl renameroo for output signals
  nios2_clock_10_out_requests_mode_select_s1 <= internal_nios2_clock_10_out_requests_mode_select_s1;
--synthesis translate_off
    --mode_select/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_0_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal nios2_clock_0_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_0_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_instruction_master_granted_nios2_clock_0_in : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_nios2_clock_0_in : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_nios2_clock_0_in : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_nios2_clock_0_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_0_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_0_in_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_clock_0_in_read : OUT STD_LOGIC;
                 signal nios2_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_0_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_0_in_write : OUT STD_LOGIC
              );
end entity nios2_clock_0_in_arbitrator;


architecture europa of nios2_clock_0_in_arbitrator is
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_nios2_clock_0_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_0_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_nios2_clock_0_in :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_nios2_clock_0_in :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_nios2_clock_0_in :  STD_LOGIC;
                signal internal_nios2_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_0_in_allgrants :  STD_LOGIC;
                signal nios2_clock_0_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_0_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_0_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_0_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_0_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_0_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_0_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_0_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_0_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_0_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_0_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_0_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_0_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_0_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_0_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_0_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_0_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_0_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_0_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_0_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_0_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_0_in_waits_for_write :  STD_LOGIC;
                signal wait_for_nios2_clock_0_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_0_in_end_xfer;
    end if;

  end process;

  nios2_clock_0_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_instruction_master_qualified_request_nios2_clock_0_in);
  --assign nios2_clock_0_in_readdata_from_sa = nios2_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_0_in_readdata_from_sa <= nios2_clock_0_in_readdata;
  internal_cpu_0_instruction_master_requests_nios2_clock_0_in <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(24 DOWNTO 15) & std_logic_vector'("000000000000000")) = std_logic_vector'("1000000001000000000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --assign nios2_clock_0_in_waitrequest_from_sa = nios2_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_0_in_waitrequest_from_sa <= nios2_clock_0_in_waitrequest;
  --nios2_clock_0_in_arb_share_counter set values, which is an e_mux
  nios2_clock_0_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_0_in_non_bursting_master_requests <= internal_cpu_0_instruction_master_requests_nios2_clock_0_in;
  --nios2_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_0_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_0_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_0_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_0_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_0_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_0_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_0_in_allgrants all slave grants, which is an e_mux
  nios2_clock_0_in_allgrants <= nios2_clock_0_in_grant_vector;
  --nios2_clock_0_in_end_xfer assignment, which is an e_assign
  nios2_clock_0_in_end_xfer <= NOT ((nios2_clock_0_in_waits_for_read OR nios2_clock_0_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_0_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_0_in <= nios2_clock_0_in_end_xfer AND (((NOT nios2_clock_0_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_0_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_0_in AND nios2_clock_0_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_0_in AND NOT nios2_clock_0_in_non_bursting_master_requests));
  --nios2_clock_0_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_0_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_0_in_arb_counter_enable) = '1' then 
        nios2_clock_0_in_arb_share_counter <= nios2_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_0_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_0_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_0_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_0_in AND NOT nios2_clock_0_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_0_in_slavearbiterlockenable <= or_reduce(nios2_clock_0_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/instruction_master nios2_clock_0/in arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= nios2_clock_0_in_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --nios2_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_0_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_0_in_arb_share_counter_next_value);
  --cpu_0/instruction_master nios2_clock_0/in arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= nios2_clock_0_in_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --nios2_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_0_in_any_continuerequest <= std_logic'('1');
  --cpu_0_instruction_master_continuerequest continued request, which is an e_assign
  cpu_0_instruction_master_continuerequest <= std_logic'('1');
  internal_cpu_0_instruction_master_qualified_request_nios2_clock_0_in <= internal_cpu_0_instruction_master_requests_nios2_clock_0_in AND NOT ((cpu_0_instruction_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_instruction_master_read_data_valid_nios2_clock_0_in, which is an e_mux
  cpu_0_instruction_master_read_data_valid_nios2_clock_0_in <= (internal_cpu_0_instruction_master_granted_nios2_clock_0_in AND cpu_0_instruction_master_read) AND NOT nios2_clock_0_in_waits_for_read;
  --assign nios2_clock_0_in_endofpacket_from_sa = nios2_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_0_in_endofpacket_from_sa <= nios2_clock_0_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_instruction_master_granted_nios2_clock_0_in <= internal_cpu_0_instruction_master_qualified_request_nios2_clock_0_in;
  --cpu_0/instruction_master saved-grant nios2_clock_0/in, which is an e_assign
  cpu_0_instruction_master_saved_grant_nios2_clock_0_in <= internal_cpu_0_instruction_master_requests_nios2_clock_0_in;
  --allow new arb cycle for nios2_clock_0/in, which is an e_assign
  nios2_clock_0_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_0_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_0_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_0_in_reset_n assignment, which is an e_assign
  nios2_clock_0_in_reset_n <= reset_n;
  --nios2_clock_0_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_0_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_0_in_begins_xfer) = '1'), nios2_clock_0_in_unreg_firsttransfer, nios2_clock_0_in_reg_firsttransfer);
  --nios2_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_0_in_unreg_firsttransfer <= NOT ((nios2_clock_0_in_slavearbiterlockenable AND nios2_clock_0_in_any_continuerequest));
  --nios2_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_0_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_0_in_begins_xfer) = '1' then 
        nios2_clock_0_in_reg_firsttransfer <= nios2_clock_0_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_0_in_beginbursttransfer_internal <= nios2_clock_0_in_begins_xfer;
  --nios2_clock_0_in_read assignment, which is an e_mux
  nios2_clock_0_in_read <= internal_cpu_0_instruction_master_granted_nios2_clock_0_in AND cpu_0_instruction_master_read;
  --nios2_clock_0_in_write assignment, which is an e_mux
  nios2_clock_0_in_write <= std_logic'('0');
  --nios2_clock_0_in_address mux, which is an e_mux
  nios2_clock_0_in_address <= cpu_0_instruction_master_address_to_slave (14 DOWNTO 0);
  --slaveid nios2_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_0_in_nativeaddress <= A_EXT (A_SRL(cpu_0_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 13);
  --d1_nios2_clock_0_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_0_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_0_in_end_xfer <= nios2_clock_0_in_end_xfer;
    end if;

  end process;

  --nios2_clock_0_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_0_in_waits_for_read <= nios2_clock_0_in_in_a_read_cycle AND internal_nios2_clock_0_in_waitrequest_from_sa;
  --nios2_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_0_in_in_a_read_cycle <= internal_cpu_0_instruction_master_granted_nios2_clock_0_in AND cpu_0_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_0_in_in_a_read_cycle;
  --nios2_clock_0_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_0_in_waits_for_write <= nios2_clock_0_in_in_a_write_cycle AND internal_nios2_clock_0_in_waitrequest_from_sa;
  --nios2_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_0_in_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_0_in_in_a_write_cycle;
  wait_for_nios2_clock_0_in_counter <= std_logic'('0');
  --nios2_clock_0_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_0_in_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 4);
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_nios2_clock_0_in <= internal_cpu_0_instruction_master_granted_nios2_clock_0_in;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_nios2_clock_0_in <= internal_cpu_0_instruction_master_qualified_request_nios2_clock_0_in;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_nios2_clock_0_in <= internal_cpu_0_instruction_master_requests_nios2_clock_0_in;
  --vhdl renameroo for output signals
  nios2_clock_0_in_waitrequest_from_sa <= internal_nios2_clock_0_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_0/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_0_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_onchip_mem_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_0_out_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_0_out_granted_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_0_out_qualified_request_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_0_out_read : IN STD_LOGIC;
                 signal nios2_clock_0_out_read_data_valid_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_0_out_requests_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_0_out_write : IN STD_LOGIC;
                 signal nios2_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal onchip_mem_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_0_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_0_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_0_out_arbitrator;


architecture europa of nios2_clock_0_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal internal_nios2_clock_0_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_0_out_address_last_time :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_0_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_0_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_0_out_run :  STD_LOGIC;
                signal nios2_clock_0_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_0_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((nios2_clock_0_out_qualified_request_onchip_mem_s1 OR nios2_clock_0_out_read_data_valid_onchip_mem_s1) OR NOT nios2_clock_0_out_requests_onchip_mem_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_0_out_granted_onchip_mem_s1 OR NOT nios2_clock_0_out_qualified_request_onchip_mem_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT nios2_clock_0_out_qualified_request_onchip_mem_s1 OR NOT nios2_clock_0_out_read) OR ((nios2_clock_0_out_read_data_valid_onchip_mem_s1 AND nios2_clock_0_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_0_out_qualified_request_onchip_mem_s1 OR NOT ((nios2_clock_0_out_read OR nios2_clock_0_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_0_out_read OR nios2_clock_0_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_0_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_0_out_address_to_slave <= nios2_clock_0_out_address;
  --nios2_clock_0/out readdata mux, which is an e_mux
  nios2_clock_0_out_readdata <= onchip_mem_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_0_out_waitrequest <= NOT nios2_clock_0_out_run;
  --nios2_clock_0_out_reset_n assignment, which is an e_assign
  nios2_clock_0_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_0_out_address_to_slave <= internal_nios2_clock_0_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_0_out_waitrequest <= internal_nios2_clock_0_out_waitrequest;
--synthesis translate_off
    --nios2_clock_0_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_0_out_address_last_time <= std_logic_vector'("000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_0_out_address_last_time <= nios2_clock_0_out_address;
      end if;

    end process;

    --nios2_clock_0/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_0_out_waitrequest AND ((nios2_clock_0_out_read OR nios2_clock_0_out_write));
      end if;

    end process;

    --nios2_clock_0_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_0_out_address /= nios2_clock_0_out_address_last_time))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("nios2_clock_0_out_address did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_0_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_0_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_0_out_byteenable_last_time <= nios2_clock_0_out_byteenable;
      end if;

    end process;

    --nios2_clock_0_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_0_out_byteenable /= nios2_clock_0_out_byteenable_last_time))))) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("nios2_clock_0_out_byteenable did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_0_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_0_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_0_out_read_last_time <= nios2_clock_0_out_read;
      end if;

    end process;

    --nios2_clock_0_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_0_out_read) /= std_logic'(nios2_clock_0_out_read_last_time)))))) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("nios2_clock_0_out_read did not heed wait!!!"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_0_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_0_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_0_out_write_last_time <= nios2_clock_0_out_write;
      end if;

    end process;

    --nios2_clock_0_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_0_out_write) /= std_logic'(nios2_clock_0_out_write_last_time)))))) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("nios2_clock_0_out_write did not heed wait!!!"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_0_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_0_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_0_out_writedata_last_time <= nios2_clock_0_out_writedata;
      end if;

    end process;

    --nios2_clock_0_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_0_out_writedata /= nios2_clock_0_out_writedata_last_time)))) AND nios2_clock_0_out_write)) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("nios2_clock_0_out_writedata did not heed wait!!!"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_1_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_1_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_1_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_1_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_1_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_1_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_1_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_1_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_1_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_1_in_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_1_in_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_clock_1_in_read : OUT STD_LOGIC;
                 signal nios2_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_1_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_1_in_write : OUT STD_LOGIC;
                 signal nios2_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_clock_1_in_arbitrator;


architecture europa of nios2_clock_1_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_1_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_1_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_1_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_1_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_1_in :  STD_LOGIC;
                signal internal_nios2_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_1_in_allgrants :  STD_LOGIC;
                signal nios2_clock_1_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_1_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_1_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_1_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_1_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_1_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_1_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_1_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_1_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_1_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_1_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_1_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_1_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_1_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_1_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_1_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_1_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_1_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_1_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_1_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_1_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_1_in_waits_for_write :  STD_LOGIC;
                signal wait_for_nios2_clock_1_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_1_in_end_xfer;
    end if;

  end process;

  nios2_clock_1_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_1_in);
  --assign nios2_clock_1_in_readdata_from_sa = nios2_clock_1_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_1_in_readdata_from_sa <= nios2_clock_1_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_1_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 15) & std_logic_vector'("000000000000000")) = std_logic_vector'("1000000001000000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_1_in_waitrequest_from_sa = nios2_clock_1_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_1_in_waitrequest_from_sa <= nios2_clock_1_in_waitrequest;
  --nios2_clock_1_in_arb_share_counter set values, which is an e_mux
  nios2_clock_1_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_1_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_1_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_1_in;
  --nios2_clock_1_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_1_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_1_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_1_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_1_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_1_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_1_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_1_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_1_in_allgrants all slave grants, which is an e_mux
  nios2_clock_1_in_allgrants <= nios2_clock_1_in_grant_vector;
  --nios2_clock_1_in_end_xfer assignment, which is an e_assign
  nios2_clock_1_in_end_xfer <= NOT ((nios2_clock_1_in_waits_for_read OR nios2_clock_1_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_1_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_1_in <= nios2_clock_1_in_end_xfer AND (((NOT nios2_clock_1_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_1_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_1_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_1_in AND nios2_clock_1_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_1_in AND NOT nios2_clock_1_in_non_bursting_master_requests));
  --nios2_clock_1_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_1_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_1_in_arb_counter_enable) = '1' then 
        nios2_clock_1_in_arb_share_counter <= nios2_clock_1_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_1_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_1_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_1_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_1_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_1_in AND NOT nios2_clock_1_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_1_in_slavearbiterlockenable <= or_reduce(nios2_clock_1_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_1/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_1_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_1_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_1_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_1_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_1/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_1_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_1_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_1_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_1_in <= internal_cpu_0_data_master_requests_nios2_clock_1_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_1_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_1_in <= (internal_cpu_0_data_master_granted_nios2_clock_1_in AND cpu_0_data_master_read) AND NOT nios2_clock_1_in_waits_for_read;
  --nios2_clock_1_in_writedata mux, which is an e_mux
  nios2_clock_1_in_writedata <= cpu_0_data_master_writedata;
  --assign nios2_clock_1_in_endofpacket_from_sa = nios2_clock_1_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_1_in_endofpacket_from_sa <= nios2_clock_1_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_1_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_1_in;
  --cpu_0/data_master saved-grant nios2_clock_1/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_1_in <= internal_cpu_0_data_master_requests_nios2_clock_1_in;
  --allow new arb cycle for nios2_clock_1/in, which is an e_assign
  nios2_clock_1_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_1_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_1_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_1_in_reset_n assignment, which is an e_assign
  nios2_clock_1_in_reset_n <= reset_n;
  --nios2_clock_1_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_1_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_1_in_begins_xfer) = '1'), nios2_clock_1_in_unreg_firsttransfer, nios2_clock_1_in_reg_firsttransfer);
  --nios2_clock_1_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_1_in_unreg_firsttransfer <= NOT ((nios2_clock_1_in_slavearbiterlockenable AND nios2_clock_1_in_any_continuerequest));
  --nios2_clock_1_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_1_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_1_in_begins_xfer) = '1' then 
        nios2_clock_1_in_reg_firsttransfer <= nios2_clock_1_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_1_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_1_in_beginbursttransfer_internal <= nios2_clock_1_in_begins_xfer;
  --nios2_clock_1_in_read assignment, which is an e_mux
  nios2_clock_1_in_read <= internal_cpu_0_data_master_granted_nios2_clock_1_in AND cpu_0_data_master_read;
  --nios2_clock_1_in_write assignment, which is an e_mux
  nios2_clock_1_in_write <= internal_cpu_0_data_master_granted_nios2_clock_1_in AND cpu_0_data_master_write;
  --nios2_clock_1_in_address mux, which is an e_mux
  nios2_clock_1_in_address <= cpu_0_data_master_address_to_slave (14 DOWNTO 0);
  --slaveid nios2_clock_1_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_1_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 13);
  --d1_nios2_clock_1_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_1_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_1_in_end_xfer <= nios2_clock_1_in_end_xfer;
    end if;

  end process;

  --nios2_clock_1_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_1_in_waits_for_read <= nios2_clock_1_in_in_a_read_cycle AND internal_nios2_clock_1_in_waitrequest_from_sa;
  --nios2_clock_1_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_1_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_1_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_1_in_in_a_read_cycle;
  --nios2_clock_1_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_1_in_waits_for_write <= nios2_clock_1_in_in_a_write_cycle AND internal_nios2_clock_1_in_waitrequest_from_sa;
  --nios2_clock_1_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_1_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_1_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_1_in_in_a_write_cycle;
  wait_for_nios2_clock_1_in_counter <= std_logic'('0');
  --nios2_clock_1_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_1_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_1_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_1_in <= internal_cpu_0_data_master_granted_nios2_clock_1_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_1_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_1_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_1_in <= internal_cpu_0_data_master_requests_nios2_clock_1_in;
  --vhdl renameroo for output signals
  nios2_clock_1_in_waitrequest_from_sa <= internal_nios2_clock_1_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_1/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_1_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_onchip_mem_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_1_out_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_1_out_granted_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_1_out_qualified_request_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_1_out_read : IN STD_LOGIC;
                 signal nios2_clock_1_out_read_data_valid_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_1_out_requests_onchip_mem_s1 : IN STD_LOGIC;
                 signal nios2_clock_1_out_write : IN STD_LOGIC;
                 signal nios2_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal onchip_mem_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_1_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_1_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_1_out_arbitrator;


architecture europa of nios2_clock_1_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal internal_nios2_clock_1_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_1_out_address_last_time :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_1_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_1_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_1_out_run :  STD_LOGIC;
                signal nios2_clock_1_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_1_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((nios2_clock_1_out_qualified_request_onchip_mem_s1 OR nios2_clock_1_out_read_data_valid_onchip_mem_s1) OR NOT nios2_clock_1_out_requests_onchip_mem_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_1_out_granted_onchip_mem_s1 OR NOT nios2_clock_1_out_qualified_request_onchip_mem_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT nios2_clock_1_out_qualified_request_onchip_mem_s1 OR NOT nios2_clock_1_out_read) OR ((nios2_clock_1_out_read_data_valid_onchip_mem_s1 AND nios2_clock_1_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_1_out_qualified_request_onchip_mem_s1 OR NOT ((nios2_clock_1_out_read OR nios2_clock_1_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_1_out_read OR nios2_clock_1_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_1_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_1_out_address_to_slave <= nios2_clock_1_out_address;
  --nios2_clock_1/out readdata mux, which is an e_mux
  nios2_clock_1_out_readdata <= onchip_mem_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_1_out_waitrequest <= NOT nios2_clock_1_out_run;
  --nios2_clock_1_out_reset_n assignment, which is an e_assign
  nios2_clock_1_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_1_out_address_to_slave <= internal_nios2_clock_1_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_1_out_waitrequest <= internal_nios2_clock_1_out_waitrequest;
--synthesis translate_off
    --nios2_clock_1_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_1_out_address_last_time <= std_logic_vector'("000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_1_out_address_last_time <= nios2_clock_1_out_address;
      end if;

    end process;

    --nios2_clock_1/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_1_out_waitrequest AND ((nios2_clock_1_out_read OR nios2_clock_1_out_write));
      end if;

    end process;

    --nios2_clock_1_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_1_out_address /= nios2_clock_1_out_address_last_time))))) = '1' then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("nios2_clock_1_out_address did not heed wait!!!"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_1_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_1_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_1_out_byteenable_last_time <= nios2_clock_1_out_byteenable;
      end if;

    end process;

    --nios2_clock_1_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_1_out_byteenable /= nios2_clock_1_out_byteenable_last_time))))) = '1' then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("nios2_clock_1_out_byteenable did not heed wait!!!"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_1_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_1_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_1_out_read_last_time <= nios2_clock_1_out_read;
      end if;

    end process;

    --nios2_clock_1_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_1_out_read) /= std_logic'(nios2_clock_1_out_read_last_time)))))) = '1' then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("nios2_clock_1_out_read did not heed wait!!!"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_1_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_1_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_1_out_write_last_time <= nios2_clock_1_out_write;
      end if;

    end process;

    --nios2_clock_1_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_1_out_write) /= std_logic'(nios2_clock_1_out_write_last_time)))))) = '1' then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("nios2_clock_1_out_write did not heed wait!!!"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_1_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_1_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_1_out_writedata_last_time <= nios2_clock_1_out_writedata;
      end if;

    end process;

    --nios2_clock_1_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_1_out_writedata /= nios2_clock_1_out_writedata_last_time)))) AND nios2_clock_1_out_write)) = '1' then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("nios2_clock_1_out_writedata did not heed wait!!!"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_10_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_10_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_10_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_10_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_10_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_10_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_10_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_10_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_10_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_10_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_10_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_in_read : OUT STD_LOGIC;
                 signal nios2_clock_10_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_10_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_10_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_10_in_write : OUT STD_LOGIC;
                 signal nios2_clock_10_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios2_clock_10_in_arbitrator;


architecture europa of nios2_clock_10_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_10_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_10_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_10_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_10_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_10_in :  STD_LOGIC;
                signal internal_nios2_clock_10_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_10_in_allgrants :  STD_LOGIC;
                signal nios2_clock_10_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_10_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_10_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_10_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_10_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_10_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_10_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_10_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_10_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_10_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_10_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_10_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_10_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_10_in_pretend_byte_enable :  STD_LOGIC;
                signal nios2_clock_10_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_10_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_10_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_10_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_10_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_10_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_10_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_10_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_10_in_end_xfer;
    end if;

  end process;

  nios2_clock_10_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_10_in);
  --assign nios2_clock_10_in_readdata_from_sa = nios2_clock_10_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_10_in_readdata_from_sa <= nios2_clock_10_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_10_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000001010000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_10_in_waitrequest_from_sa = nios2_clock_10_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_10_in_waitrequest_from_sa <= nios2_clock_10_in_waitrequest;
  --nios2_clock_10_in_arb_share_counter set values, which is an e_mux
  nios2_clock_10_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_10_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_10_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_10_in;
  --nios2_clock_10_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_10_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_10_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_10_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_10_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_10_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_10_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_10_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_10_in_allgrants all slave grants, which is an e_mux
  nios2_clock_10_in_allgrants <= nios2_clock_10_in_grant_vector;
  --nios2_clock_10_in_end_xfer assignment, which is an e_assign
  nios2_clock_10_in_end_xfer <= NOT ((nios2_clock_10_in_waits_for_read OR nios2_clock_10_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_10_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_10_in <= nios2_clock_10_in_end_xfer AND (((NOT nios2_clock_10_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_10_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_10_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_10_in AND nios2_clock_10_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_10_in AND NOT nios2_clock_10_in_non_bursting_master_requests));
  --nios2_clock_10_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_10_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_10_in_arb_counter_enable) = '1' then 
        nios2_clock_10_in_arb_share_counter <= nios2_clock_10_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_10_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_10_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_10_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_10_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_10_in AND NOT nios2_clock_10_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_10_in_slavearbiterlockenable <= or_reduce(nios2_clock_10_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_10/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_10_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_10_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_10_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_10_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_10/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_10_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_10_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_10_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_10_in <= internal_cpu_0_data_master_requests_nios2_clock_10_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_10_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_10_in <= (internal_cpu_0_data_master_granted_nios2_clock_10_in AND cpu_0_data_master_read) AND NOT nios2_clock_10_in_waits_for_read;
  --nios2_clock_10_in_writedata mux, which is an e_mux
  nios2_clock_10_in_writedata <= cpu_0_data_master_writedata (7 DOWNTO 0);
  --assign nios2_clock_10_in_endofpacket_from_sa = nios2_clock_10_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_10_in_endofpacket_from_sa <= nios2_clock_10_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_10_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_10_in;
  --cpu_0/data_master saved-grant nios2_clock_10/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_10_in <= internal_cpu_0_data_master_requests_nios2_clock_10_in;
  --allow new arb cycle for nios2_clock_10/in, which is an e_assign
  nios2_clock_10_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_10_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_10_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_10_in_reset_n assignment, which is an e_assign
  nios2_clock_10_in_reset_n <= reset_n;
  --nios2_clock_10_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_10_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_10_in_begins_xfer) = '1'), nios2_clock_10_in_unreg_firsttransfer, nios2_clock_10_in_reg_firsttransfer);
  --nios2_clock_10_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_10_in_unreg_firsttransfer <= NOT ((nios2_clock_10_in_slavearbiterlockenable AND nios2_clock_10_in_any_continuerequest));
  --nios2_clock_10_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_10_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_10_in_begins_xfer) = '1' then 
        nios2_clock_10_in_reg_firsttransfer <= nios2_clock_10_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_10_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_10_in_beginbursttransfer_internal <= nios2_clock_10_in_begins_xfer;
  --nios2_clock_10_in_read assignment, which is an e_mux
  nios2_clock_10_in_read <= internal_cpu_0_data_master_granted_nios2_clock_10_in AND cpu_0_data_master_read;
  --nios2_clock_10_in_write assignment, which is an e_mux
  nios2_clock_10_in_write <= ((internal_cpu_0_data_master_granted_nios2_clock_10_in AND cpu_0_data_master_write)) AND nios2_clock_10_in_pretend_byte_enable;
  shifted_address_to_nios2_clock_10_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_10_in_address mux, which is an e_mux
  nios2_clock_10_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_10_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --slaveid nios2_clock_10_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_10_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_10_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_10_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_10_in_end_xfer <= nios2_clock_10_in_end_xfer;
    end if;

  end process;

  --nios2_clock_10_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_10_in_waits_for_read <= nios2_clock_10_in_in_a_read_cycle AND internal_nios2_clock_10_in_waitrequest_from_sa;
  --nios2_clock_10_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_10_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_10_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_10_in_in_a_read_cycle;
  --nios2_clock_10_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_10_in_waits_for_write <= nios2_clock_10_in_in_a_write_cycle AND internal_nios2_clock_10_in_waitrequest_from_sa;
  --nios2_clock_10_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_10_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_10_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_10_in_in_a_write_cycle;
  wait_for_nios2_clock_10_in_counter <= std_logic'('0');
  --nios2_clock_10_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios2_clock_10_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_10_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_10_in <= internal_cpu_0_data_master_granted_nios2_clock_10_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_10_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_10_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_10_in <= internal_cpu_0_data_master_requests_nios2_clock_10_in;
  --vhdl renameroo for output signals
  nios2_clock_10_in_waitrequest_from_sa <= internal_nios2_clock_10_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_10/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_10_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_mode_select_s1_end_xfer : IN STD_LOGIC;
                 signal mode_select_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_out_granted_mode_select_s1 : IN STD_LOGIC;
                 signal nios2_clock_10_out_qualified_request_mode_select_s1 : IN STD_LOGIC;
                 signal nios2_clock_10_out_read : IN STD_LOGIC;
                 signal nios2_clock_10_out_read_data_valid_mode_select_s1 : IN STD_LOGIC;
                 signal nios2_clock_10_out_requests_mode_select_s1 : IN STD_LOGIC;
                 signal nios2_clock_10_out_write : IN STD_LOGIC;
                 signal nios2_clock_10_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_10_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_10_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_10_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_10_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_10_out_arbitrator;


architecture europa of nios2_clock_10_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_10_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_clock_10_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_10_out_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_10_out_run :  STD_LOGIC;
                signal nios2_clock_10_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_10_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_10_out_qualified_request_mode_select_s1 OR NOT nios2_clock_10_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_mode_select_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_10_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_10_out_qualified_request_mode_select_s1 OR NOT nios2_clock_10_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_10_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_10_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_10_out_address_to_slave <= nios2_clock_10_out_address;
  --nios2_clock_10/out readdata mux, which is an e_mux
  nios2_clock_10_out_readdata <= std_logic_vector'("000000") & (mode_select_s1_readdata_from_sa);
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_10_out_waitrequest <= NOT nios2_clock_10_out_run;
  --nios2_clock_10_out_reset_n assignment, which is an e_assign
  nios2_clock_10_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_10_out_address_to_slave <= internal_nios2_clock_10_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_10_out_waitrequest <= internal_nios2_clock_10_out_waitrequest;
--synthesis translate_off
    --nios2_clock_10_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_10_out_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_10_out_address_last_time <= nios2_clock_10_out_address;
      end if;

    end process;

    --nios2_clock_10/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_10_out_waitrequest AND ((nios2_clock_10_out_read OR nios2_clock_10_out_write));
      end if;

    end process;

    --nios2_clock_10_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_10_out_address /= nios2_clock_10_out_address_last_time))))) = '1' then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("nios2_clock_10_out_address did not heed wait!!!"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_10_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_10_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_10_out_read_last_time <= nios2_clock_10_out_read;
      end if;

    end process;

    --nios2_clock_10_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_10_out_read) /= std_logic'(nios2_clock_10_out_read_last_time)))))) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("nios2_clock_10_out_read did not heed wait!!!"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_10_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_10_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_10_out_write_last_time <= nios2_clock_10_out_write;
      end if;

    end process;

    --nios2_clock_10_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_10_out_write) /= std_logic'(nios2_clock_10_out_write_last_time)))))) = '1' then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("nios2_clock_10_out_write did not heed wait!!!"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_10_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_10_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios2_clock_10_out_writedata_last_time <= nios2_clock_10_out_writedata;
      end if;

    end process;

    --nios2_clock_10_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_10_out_writedata /= nios2_clock_10_out_writedata_last_time)))) AND nios2_clock_10_out_write)) = '1' then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("nios2_clock_10_out_writedata did not heed wait!!!"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_11_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_11_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_11_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_11_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_11_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_11_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_11_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_11_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_11_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_11_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_11_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_11_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_11_in_read : OUT STD_LOGIC;
                 signal nios2_clock_11_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_11_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_11_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_11_in_write : OUT STD_LOGIC;
                 signal nios2_clock_11_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios2_clock_11_in_arbitrator;


architecture europa of nios2_clock_11_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_11_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_11_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_11_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_11_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_11_in :  STD_LOGIC;
                signal internal_nios2_clock_11_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_11_in_allgrants :  STD_LOGIC;
                signal nios2_clock_11_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_11_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_11_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_11_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_11_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_11_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_11_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_11_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_11_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_11_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_11_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_11_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_11_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_11_in_pretend_byte_enable :  STD_LOGIC;
                signal nios2_clock_11_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_11_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_11_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_11_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_11_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_11_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_11_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_11_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_11_in_end_xfer;
    end if;

  end process;

  nios2_clock_11_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_11_in);
  --assign nios2_clock_11_in_readdata_from_sa = nios2_clock_11_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_11_in_readdata_from_sa <= nios2_clock_11_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_11_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000001100000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_11_in_waitrequest_from_sa = nios2_clock_11_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_11_in_waitrequest_from_sa <= nios2_clock_11_in_waitrequest;
  --nios2_clock_11_in_arb_share_counter set values, which is an e_mux
  nios2_clock_11_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_11_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_11_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_11_in;
  --nios2_clock_11_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_11_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_11_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_11_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_11_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_11_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_11_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_11_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_11_in_allgrants all slave grants, which is an e_mux
  nios2_clock_11_in_allgrants <= nios2_clock_11_in_grant_vector;
  --nios2_clock_11_in_end_xfer assignment, which is an e_assign
  nios2_clock_11_in_end_xfer <= NOT ((nios2_clock_11_in_waits_for_read OR nios2_clock_11_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_11_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_11_in <= nios2_clock_11_in_end_xfer AND (((NOT nios2_clock_11_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_11_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_11_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_11_in AND nios2_clock_11_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_11_in AND NOT nios2_clock_11_in_non_bursting_master_requests));
  --nios2_clock_11_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_11_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_11_in_arb_counter_enable) = '1' then 
        nios2_clock_11_in_arb_share_counter <= nios2_clock_11_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_11_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_11_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_11_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_11_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_11_in AND NOT nios2_clock_11_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_11_in_slavearbiterlockenable <= or_reduce(nios2_clock_11_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_11/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_11_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_11_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_11_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_11_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_11/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_11_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_11_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_11_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_11_in <= internal_cpu_0_data_master_requests_nios2_clock_11_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_11_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_11_in <= (internal_cpu_0_data_master_granted_nios2_clock_11_in AND cpu_0_data_master_read) AND NOT nios2_clock_11_in_waits_for_read;
  --nios2_clock_11_in_writedata mux, which is an e_mux
  nios2_clock_11_in_writedata <= cpu_0_data_master_writedata (7 DOWNTO 0);
  --assign nios2_clock_11_in_endofpacket_from_sa = nios2_clock_11_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_11_in_endofpacket_from_sa <= nios2_clock_11_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_11_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_11_in;
  --cpu_0/data_master saved-grant nios2_clock_11/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_11_in <= internal_cpu_0_data_master_requests_nios2_clock_11_in;
  --allow new arb cycle for nios2_clock_11/in, which is an e_assign
  nios2_clock_11_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_11_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_11_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_11_in_reset_n assignment, which is an e_assign
  nios2_clock_11_in_reset_n <= reset_n;
  --nios2_clock_11_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_11_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_11_in_begins_xfer) = '1'), nios2_clock_11_in_unreg_firsttransfer, nios2_clock_11_in_reg_firsttransfer);
  --nios2_clock_11_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_11_in_unreg_firsttransfer <= NOT ((nios2_clock_11_in_slavearbiterlockenable AND nios2_clock_11_in_any_continuerequest));
  --nios2_clock_11_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_11_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_11_in_begins_xfer) = '1' then 
        nios2_clock_11_in_reg_firsttransfer <= nios2_clock_11_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_11_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_11_in_beginbursttransfer_internal <= nios2_clock_11_in_begins_xfer;
  --nios2_clock_11_in_read assignment, which is an e_mux
  nios2_clock_11_in_read <= internal_cpu_0_data_master_granted_nios2_clock_11_in AND cpu_0_data_master_read;
  --nios2_clock_11_in_write assignment, which is an e_mux
  nios2_clock_11_in_write <= ((internal_cpu_0_data_master_granted_nios2_clock_11_in AND cpu_0_data_master_write)) AND nios2_clock_11_in_pretend_byte_enable;
  shifted_address_to_nios2_clock_11_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_11_in_address mux, which is an e_mux
  nios2_clock_11_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_11_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --slaveid nios2_clock_11_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_11_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_11_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_11_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_11_in_end_xfer <= nios2_clock_11_in_end_xfer;
    end if;

  end process;

  --nios2_clock_11_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_11_in_waits_for_read <= nios2_clock_11_in_in_a_read_cycle AND internal_nios2_clock_11_in_waitrequest_from_sa;
  --nios2_clock_11_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_11_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_11_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_11_in_in_a_read_cycle;
  --nios2_clock_11_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_11_in_waits_for_write <= nios2_clock_11_in_in_a_write_cycle AND internal_nios2_clock_11_in_waitrequest_from_sa;
  --nios2_clock_11_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_11_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_11_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_11_in_in_a_write_cycle;
  wait_for_nios2_clock_11_in_counter <= std_logic'('0');
  --nios2_clock_11_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios2_clock_11_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_11_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_11_in <= internal_cpu_0_data_master_granted_nios2_clock_11_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_11_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_11_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_11_in <= internal_cpu_0_data_master_requests_nios2_clock_11_in;
  --vhdl renameroo for output signals
  nios2_clock_11_in_waitrequest_from_sa <= internal_nios2_clock_11_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_11/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_11_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal comparator_pio_s1_readdata_from_sa : IN STD_LOGIC;
                 signal d1_comparator_pio_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_11_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_11_out_granted_comparator_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_11_out_qualified_request_comparator_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_11_out_read : IN STD_LOGIC;
                 signal nios2_clock_11_out_read_data_valid_comparator_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_11_out_requests_comparator_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_11_out_write : IN STD_LOGIC;
                 signal nios2_clock_11_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_11_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_11_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_11_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_11_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_11_out_arbitrator;


architecture europa of nios2_clock_11_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_11_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_clock_11_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_11_out_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_11_out_run :  STD_LOGIC;
                signal nios2_clock_11_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_11_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_11_out_qualified_request_comparator_pio_s1 OR NOT nios2_clock_11_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_comparator_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_11_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_11_out_qualified_request_comparator_pio_s1 OR NOT nios2_clock_11_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_11_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_11_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_11_out_address_to_slave <= nios2_clock_11_out_address;
  --nios2_clock_11/out readdata mux, which is an e_mux
  nios2_clock_11_out_readdata <= std_logic_vector'("0000000") & (A_TOSTDLOGICVECTOR(comparator_pio_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_11_out_waitrequest <= NOT nios2_clock_11_out_run;
  --nios2_clock_11_out_reset_n assignment, which is an e_assign
  nios2_clock_11_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_11_out_address_to_slave <= internal_nios2_clock_11_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_11_out_waitrequest <= internal_nios2_clock_11_out_waitrequest;
--synthesis translate_off
    --nios2_clock_11_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_11_out_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_11_out_address_last_time <= nios2_clock_11_out_address;
      end if;

    end process;

    --nios2_clock_11/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_11_out_waitrequest AND ((nios2_clock_11_out_read OR nios2_clock_11_out_write));
      end if;

    end process;

    --nios2_clock_11_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_11_out_address /= nios2_clock_11_out_address_last_time))))) = '1' then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("nios2_clock_11_out_address did not heed wait!!!"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_11_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_11_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_11_out_read_last_time <= nios2_clock_11_out_read;
      end if;

    end process;

    --nios2_clock_11_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_11_out_read) /= std_logic'(nios2_clock_11_out_read_last_time)))))) = '1' then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("nios2_clock_11_out_read did not heed wait!!!"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_11_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_11_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_11_out_write_last_time <= nios2_clock_11_out_write;
      end if;

    end process;

    --nios2_clock_11_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_11_out_write) /= std_logic'(nios2_clock_11_out_write_last_time)))))) = '1' then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("nios2_clock_11_out_write did not heed wait!!!"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_11_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_11_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios2_clock_11_out_writedata_last_time <= nios2_clock_11_out_writedata;
      end if;

    end process;

    --nios2_clock_11_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_11_out_writedata /= nios2_clock_11_out_writedata_last_time)))) AND nios2_clock_11_out_write)) = '1' then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("nios2_clock_11_out_writedata did not heed wait!!!"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_12_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_12_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_12_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_12_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_12_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_12_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_12_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_12_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_12_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_12_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_12_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_12_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_12_in_read : OUT STD_LOGIC;
                 signal nios2_clock_12_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_12_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_12_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_12_in_write : OUT STD_LOGIC;
                 signal nios2_clock_12_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios2_clock_12_in_arbitrator;


architecture europa of nios2_clock_12_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_12_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_12_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_12_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_12_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_12_in :  STD_LOGIC;
                signal internal_nios2_clock_12_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_12_in_allgrants :  STD_LOGIC;
                signal nios2_clock_12_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_12_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_12_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_12_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_12_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_12_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_12_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_12_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_12_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_12_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_12_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_12_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_12_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_12_in_pretend_byte_enable :  STD_LOGIC;
                signal nios2_clock_12_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_12_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_12_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_12_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_12_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_12_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_12_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_12_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_12_in_end_xfer;
    end if;

  end process;

  nios2_clock_12_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_12_in);
  --assign nios2_clock_12_in_readdata_from_sa = nios2_clock_12_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_12_in_readdata_from_sa <= nios2_clock_12_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_12_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000001110000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_12_in_waitrequest_from_sa = nios2_clock_12_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_12_in_waitrequest_from_sa <= nios2_clock_12_in_waitrequest;
  --nios2_clock_12_in_arb_share_counter set values, which is an e_mux
  nios2_clock_12_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_12_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_12_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_12_in;
  --nios2_clock_12_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_12_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_12_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_12_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_12_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_12_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_12_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_12_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_12_in_allgrants all slave grants, which is an e_mux
  nios2_clock_12_in_allgrants <= nios2_clock_12_in_grant_vector;
  --nios2_clock_12_in_end_xfer assignment, which is an e_assign
  nios2_clock_12_in_end_xfer <= NOT ((nios2_clock_12_in_waits_for_read OR nios2_clock_12_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_12_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_12_in <= nios2_clock_12_in_end_xfer AND (((NOT nios2_clock_12_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_12_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_12_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_12_in AND nios2_clock_12_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_12_in AND NOT nios2_clock_12_in_non_bursting_master_requests));
  --nios2_clock_12_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_12_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_12_in_arb_counter_enable) = '1' then 
        nios2_clock_12_in_arb_share_counter <= nios2_clock_12_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_12_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_12_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_12_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_12_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_12_in AND NOT nios2_clock_12_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_12_in_slavearbiterlockenable <= or_reduce(nios2_clock_12_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_12/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_12_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_12_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_12_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_12_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_12/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_12_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_12_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_12_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_12_in <= internal_cpu_0_data_master_requests_nios2_clock_12_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_12_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_12_in <= (internal_cpu_0_data_master_granted_nios2_clock_12_in AND cpu_0_data_master_read) AND NOT nios2_clock_12_in_waits_for_read;
  --nios2_clock_12_in_writedata mux, which is an e_mux
  nios2_clock_12_in_writedata <= cpu_0_data_master_writedata (7 DOWNTO 0);
  --assign nios2_clock_12_in_endofpacket_from_sa = nios2_clock_12_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_12_in_endofpacket_from_sa <= nios2_clock_12_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_12_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_12_in;
  --cpu_0/data_master saved-grant nios2_clock_12/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_12_in <= internal_cpu_0_data_master_requests_nios2_clock_12_in;
  --allow new arb cycle for nios2_clock_12/in, which is an e_assign
  nios2_clock_12_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_12_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_12_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_12_in_reset_n assignment, which is an e_assign
  nios2_clock_12_in_reset_n <= reset_n;
  --nios2_clock_12_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_12_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_12_in_begins_xfer) = '1'), nios2_clock_12_in_unreg_firsttransfer, nios2_clock_12_in_reg_firsttransfer);
  --nios2_clock_12_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_12_in_unreg_firsttransfer <= NOT ((nios2_clock_12_in_slavearbiterlockenable AND nios2_clock_12_in_any_continuerequest));
  --nios2_clock_12_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_12_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_12_in_begins_xfer) = '1' then 
        nios2_clock_12_in_reg_firsttransfer <= nios2_clock_12_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_12_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_12_in_beginbursttransfer_internal <= nios2_clock_12_in_begins_xfer;
  --nios2_clock_12_in_read assignment, which is an e_mux
  nios2_clock_12_in_read <= internal_cpu_0_data_master_granted_nios2_clock_12_in AND cpu_0_data_master_read;
  --nios2_clock_12_in_write assignment, which is an e_mux
  nios2_clock_12_in_write <= ((internal_cpu_0_data_master_granted_nios2_clock_12_in AND cpu_0_data_master_write)) AND nios2_clock_12_in_pretend_byte_enable;
  shifted_address_to_nios2_clock_12_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_12_in_address mux, which is an e_mux
  nios2_clock_12_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_12_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --slaveid nios2_clock_12_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_12_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_12_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_12_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_12_in_end_xfer <= nios2_clock_12_in_end_xfer;
    end if;

  end process;

  --nios2_clock_12_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_12_in_waits_for_read <= nios2_clock_12_in_in_a_read_cycle AND internal_nios2_clock_12_in_waitrequest_from_sa;
  --nios2_clock_12_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_12_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_12_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_12_in_in_a_read_cycle;
  --nios2_clock_12_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_12_in_waits_for_write <= nios2_clock_12_in_in_a_write_cycle AND internal_nios2_clock_12_in_waitrequest_from_sa;
  --nios2_clock_12_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_12_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_12_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_12_in_in_a_write_cycle;
  wait_for_nios2_clock_12_in_counter <= std_logic'('0');
  --nios2_clock_12_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios2_clock_12_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_12_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_12_in <= internal_cpu_0_data_master_granted_nios2_clock_12_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_12_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_12_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_12_in <= internal_cpu_0_data_master_requests_nios2_clock_12_in;
  --vhdl renameroo for output signals
  nios2_clock_12_in_waitrequest_from_sa <= internal_nios2_clock_12_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_12/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_12_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_12_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_12_out_granted_led_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_12_out_qualified_request_led_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_12_out_read : IN STD_LOGIC;
                 signal nios2_clock_12_out_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_12_out_requests_led_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_12_out_write : IN STD_LOGIC;
                 signal nios2_clock_12_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_12_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_12_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_12_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_12_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_12_out_arbitrator;


architecture europa of nios2_clock_12_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_12_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_clock_12_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_12_out_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_12_out_run :  STD_LOGIC;
                signal nios2_clock_12_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_12_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_12_out_qualified_request_led_pio_s1 OR NOT nios2_clock_12_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_led_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_12_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_12_out_qualified_request_led_pio_s1 OR NOT nios2_clock_12_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_12_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_12_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_12_out_address_to_slave <= nios2_clock_12_out_address;
  --nios2_clock_12/out readdata mux, which is an e_mux
  nios2_clock_12_out_readdata <= led_pio_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_12_out_waitrequest <= NOT nios2_clock_12_out_run;
  --nios2_clock_12_out_reset_n assignment, which is an e_assign
  nios2_clock_12_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_12_out_address_to_slave <= internal_nios2_clock_12_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_12_out_waitrequest <= internal_nios2_clock_12_out_waitrequest;
--synthesis translate_off
    --nios2_clock_12_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_12_out_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_12_out_address_last_time <= nios2_clock_12_out_address;
      end if;

    end process;

    --nios2_clock_12/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_12_out_waitrequest AND ((nios2_clock_12_out_read OR nios2_clock_12_out_write));
      end if;

    end process;

    --nios2_clock_12_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_12_out_address /= nios2_clock_12_out_address_last_time))))) = '1' then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("nios2_clock_12_out_address did not heed wait!!!"));
          write(output, write_line27.all);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_12_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_12_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_12_out_read_last_time <= nios2_clock_12_out_read;
      end if;

    end process;

    --nios2_clock_12_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_12_out_read) /= std_logic'(nios2_clock_12_out_read_last_time)))))) = '1' then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("nios2_clock_12_out_read did not heed wait!!!"));
          write(output, write_line28.all);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_12_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_12_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_12_out_write_last_time <= nios2_clock_12_out_write;
      end if;

    end process;

    --nios2_clock_12_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_12_out_write) /= std_logic'(nios2_clock_12_out_write_last_time)))))) = '1' then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("nios2_clock_12_out_write did not heed wait!!!"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_12_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_12_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios2_clock_12_out_writedata_last_time <= nios2_clock_12_out_writedata;
      end if;

    end process;

    --nios2_clock_12_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_12_out_writedata /= nios2_clock_12_out_writedata_last_time)))) AND nios2_clock_12_out_write)) = '1' then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("nios2_clock_12_out_writedata did not heed wait!!!"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_13_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_13_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_13_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_13_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_13_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_13_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_13_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_13_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_13_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_13_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_13_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_13_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_13_in_read : OUT STD_LOGIC;
                 signal nios2_clock_13_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_13_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_13_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_13_in_write : OUT STD_LOGIC;
                 signal nios2_clock_13_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios2_clock_13_in_arbitrator;


architecture europa of nios2_clock_13_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_13_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_13_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_13_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_13_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_13_in :  STD_LOGIC;
                signal internal_nios2_clock_13_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_13_in_allgrants :  STD_LOGIC;
                signal nios2_clock_13_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_13_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_13_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_13_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_13_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_13_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_13_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_13_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_13_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_13_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_13_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_13_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_13_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_13_in_pretend_byte_enable :  STD_LOGIC;
                signal nios2_clock_13_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_13_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_13_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_13_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_13_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_13_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_13_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_13_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_13_in_end_xfer;
    end if;

  end process;

  nios2_clock_13_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_13_in);
  --assign nios2_clock_13_in_readdata_from_sa = nios2_clock_13_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_13_in_readdata_from_sa <= nios2_clock_13_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_13_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000010000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_13_in_waitrequest_from_sa = nios2_clock_13_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_13_in_waitrequest_from_sa <= nios2_clock_13_in_waitrequest;
  --nios2_clock_13_in_arb_share_counter set values, which is an e_mux
  nios2_clock_13_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_13_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_13_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_13_in;
  --nios2_clock_13_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_13_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_13_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_13_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_13_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_13_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_13_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_13_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_13_in_allgrants all slave grants, which is an e_mux
  nios2_clock_13_in_allgrants <= nios2_clock_13_in_grant_vector;
  --nios2_clock_13_in_end_xfer assignment, which is an e_assign
  nios2_clock_13_in_end_xfer <= NOT ((nios2_clock_13_in_waits_for_read OR nios2_clock_13_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_13_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_13_in <= nios2_clock_13_in_end_xfer AND (((NOT nios2_clock_13_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_13_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_13_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_13_in AND nios2_clock_13_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_13_in AND NOT nios2_clock_13_in_non_bursting_master_requests));
  --nios2_clock_13_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_13_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_13_in_arb_counter_enable) = '1' then 
        nios2_clock_13_in_arb_share_counter <= nios2_clock_13_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_13_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_13_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_13_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_13_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_13_in AND NOT nios2_clock_13_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_13_in_slavearbiterlockenable <= or_reduce(nios2_clock_13_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_13/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_13_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_13_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_13_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_13_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_13/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_13_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_13_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_13_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_13_in <= internal_cpu_0_data_master_requests_nios2_clock_13_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_13_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_13_in <= (internal_cpu_0_data_master_granted_nios2_clock_13_in AND cpu_0_data_master_read) AND NOT nios2_clock_13_in_waits_for_read;
  --nios2_clock_13_in_writedata mux, which is an e_mux
  nios2_clock_13_in_writedata <= cpu_0_data_master_writedata (7 DOWNTO 0);
  --assign nios2_clock_13_in_endofpacket_from_sa = nios2_clock_13_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_13_in_endofpacket_from_sa <= nios2_clock_13_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_13_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_13_in;
  --cpu_0/data_master saved-grant nios2_clock_13/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_13_in <= internal_cpu_0_data_master_requests_nios2_clock_13_in;
  --allow new arb cycle for nios2_clock_13/in, which is an e_assign
  nios2_clock_13_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_13_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_13_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_13_in_reset_n assignment, which is an e_assign
  nios2_clock_13_in_reset_n <= reset_n;
  --nios2_clock_13_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_13_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_13_in_begins_xfer) = '1'), nios2_clock_13_in_unreg_firsttransfer, nios2_clock_13_in_reg_firsttransfer);
  --nios2_clock_13_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_13_in_unreg_firsttransfer <= NOT ((nios2_clock_13_in_slavearbiterlockenable AND nios2_clock_13_in_any_continuerequest));
  --nios2_clock_13_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_13_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_13_in_begins_xfer) = '1' then 
        nios2_clock_13_in_reg_firsttransfer <= nios2_clock_13_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_13_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_13_in_beginbursttransfer_internal <= nios2_clock_13_in_begins_xfer;
  --nios2_clock_13_in_read assignment, which is an e_mux
  nios2_clock_13_in_read <= internal_cpu_0_data_master_granted_nios2_clock_13_in AND cpu_0_data_master_read;
  --nios2_clock_13_in_write assignment, which is an e_mux
  nios2_clock_13_in_write <= ((internal_cpu_0_data_master_granted_nios2_clock_13_in AND cpu_0_data_master_write)) AND nios2_clock_13_in_pretend_byte_enable;
  shifted_address_to_nios2_clock_13_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_13_in_address mux, which is an e_mux
  nios2_clock_13_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_13_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --slaveid nios2_clock_13_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_13_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_13_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_13_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_13_in_end_xfer <= nios2_clock_13_in_end_xfer;
    end if;

  end process;

  --nios2_clock_13_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_13_in_waits_for_read <= nios2_clock_13_in_in_a_read_cycle AND internal_nios2_clock_13_in_waitrequest_from_sa;
  --nios2_clock_13_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_13_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_13_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_13_in_in_a_read_cycle;
  --nios2_clock_13_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_13_in_waits_for_write <= nios2_clock_13_in_in_a_write_cycle AND internal_nios2_clock_13_in_waitrequest_from_sa;
  --nios2_clock_13_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_13_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_13_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_13_in_in_a_write_cycle;
  wait_for_nios2_clock_13_in_counter <= std_logic'('0');
  --nios2_clock_13_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios2_clock_13_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_13_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_13_in <= internal_cpu_0_data_master_granted_nios2_clock_13_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_13_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_13_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_13_in <= internal_cpu_0_data_master_requests_nios2_clock_13_in;
  --vhdl renameroo for output signals
  nios2_clock_13_in_waitrequest_from_sa <= internal_nios2_clock_13_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_13/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_13_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_gen_code_strobe_s1_end_xfer : IN STD_LOGIC;
                 signal gen_code_strobe_s1_readdata_from_sa : IN STD_LOGIC;
                 signal nios2_clock_13_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_13_out_granted_gen_code_strobe_s1 : IN STD_LOGIC;
                 signal nios2_clock_13_out_qualified_request_gen_code_strobe_s1 : IN STD_LOGIC;
                 signal nios2_clock_13_out_read : IN STD_LOGIC;
                 signal nios2_clock_13_out_read_data_valid_gen_code_strobe_s1 : IN STD_LOGIC;
                 signal nios2_clock_13_out_requests_gen_code_strobe_s1 : IN STD_LOGIC;
                 signal nios2_clock_13_out_write : IN STD_LOGIC;
                 signal nios2_clock_13_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_13_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_13_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_13_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_13_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_13_out_arbitrator;


architecture europa of nios2_clock_13_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_13_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_clock_13_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_13_out_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_13_out_run :  STD_LOGIC;
                signal nios2_clock_13_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_13_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_13_out_qualified_request_gen_code_strobe_s1 OR NOT nios2_clock_13_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_gen_code_strobe_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_13_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_13_out_qualified_request_gen_code_strobe_s1 OR NOT nios2_clock_13_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_13_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_13_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_13_out_address_to_slave <= nios2_clock_13_out_address;
  --nios2_clock_13/out readdata mux, which is an e_mux
  nios2_clock_13_out_readdata <= std_logic_vector'("0000000") & (A_TOSTDLOGICVECTOR(gen_code_strobe_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_13_out_waitrequest <= NOT nios2_clock_13_out_run;
  --nios2_clock_13_out_reset_n assignment, which is an e_assign
  nios2_clock_13_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_13_out_address_to_slave <= internal_nios2_clock_13_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_13_out_waitrequest <= internal_nios2_clock_13_out_waitrequest;
--synthesis translate_off
    --nios2_clock_13_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_13_out_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_13_out_address_last_time <= nios2_clock_13_out_address;
      end if;

    end process;

    --nios2_clock_13/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_13_out_waitrequest AND ((nios2_clock_13_out_read OR nios2_clock_13_out_write));
      end if;

    end process;

    --nios2_clock_13_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_13_out_address /= nios2_clock_13_out_address_last_time))))) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("nios2_clock_13_out_address did not heed wait!!!"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_13_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_13_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_13_out_read_last_time <= nios2_clock_13_out_read;
      end if;

    end process;

    --nios2_clock_13_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_13_out_read) /= std_logic'(nios2_clock_13_out_read_last_time)))))) = '1' then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("nios2_clock_13_out_read did not heed wait!!!"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_13_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_13_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_13_out_write_last_time <= nios2_clock_13_out_write;
      end if;

    end process;

    --nios2_clock_13_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_13_out_write) /= std_logic'(nios2_clock_13_out_write_last_time)))))) = '1' then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("nios2_clock_13_out_write did not heed wait!!!"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_13_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_13_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios2_clock_13_out_writedata_last_time <= nios2_clock_13_out_writedata;
      end if;

    end process;

    --nios2_clock_13_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_13_out_writedata /= nios2_clock_13_out_writedata_last_time)))) AND nios2_clock_13_out_write)) = '1' then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("nios2_clock_13_out_writedata did not heed wait!!!"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_14_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_14_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_14_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_14_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_14_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_14_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_14_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_14_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_14_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_14_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_14_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_14_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_14_in_read : OUT STD_LOGIC;
                 signal nios2_clock_14_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_14_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_14_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_14_in_write : OUT STD_LOGIC;
                 signal nios2_clock_14_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios2_clock_14_in_arbitrator;


architecture europa of nios2_clock_14_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_14_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_14_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_14_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_14_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_14_in :  STD_LOGIC;
                signal internal_nios2_clock_14_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_14_in_allgrants :  STD_LOGIC;
                signal nios2_clock_14_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_14_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_14_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_14_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_14_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_14_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_14_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_14_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_14_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_14_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_14_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_14_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_14_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_14_in_pretend_byte_enable :  STD_LOGIC;
                signal nios2_clock_14_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_14_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_14_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_14_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_14_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_14_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_14_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_14_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_14_in_end_xfer;
    end if;

  end process;

  nios2_clock_14_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_14_in);
  --assign nios2_clock_14_in_readdata_from_sa = nios2_clock_14_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_14_in_readdata_from_sa <= nios2_clock_14_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_14_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000010010000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_14_in_waitrequest_from_sa = nios2_clock_14_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_14_in_waitrequest_from_sa <= nios2_clock_14_in_waitrequest;
  --nios2_clock_14_in_arb_share_counter set values, which is an e_mux
  nios2_clock_14_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_14_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_14_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_14_in;
  --nios2_clock_14_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_14_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_14_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_14_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_14_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_14_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_14_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_14_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_14_in_allgrants all slave grants, which is an e_mux
  nios2_clock_14_in_allgrants <= nios2_clock_14_in_grant_vector;
  --nios2_clock_14_in_end_xfer assignment, which is an e_assign
  nios2_clock_14_in_end_xfer <= NOT ((nios2_clock_14_in_waits_for_read OR nios2_clock_14_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_14_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_14_in <= nios2_clock_14_in_end_xfer AND (((NOT nios2_clock_14_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_14_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_14_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_14_in AND nios2_clock_14_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_14_in AND NOT nios2_clock_14_in_non_bursting_master_requests));
  --nios2_clock_14_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_14_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_14_in_arb_counter_enable) = '1' then 
        nios2_clock_14_in_arb_share_counter <= nios2_clock_14_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_14_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_14_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_14_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_14_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_14_in AND NOT nios2_clock_14_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_14_in_slavearbiterlockenable <= or_reduce(nios2_clock_14_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_14/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_14_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_14_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_14_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_14_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_14/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_14_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_14_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_14_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_14_in <= internal_cpu_0_data_master_requests_nios2_clock_14_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_14_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_14_in <= (internal_cpu_0_data_master_granted_nios2_clock_14_in AND cpu_0_data_master_read) AND NOT nios2_clock_14_in_waits_for_read;
  --nios2_clock_14_in_writedata mux, which is an e_mux
  nios2_clock_14_in_writedata <= cpu_0_data_master_writedata (7 DOWNTO 0);
  --assign nios2_clock_14_in_endofpacket_from_sa = nios2_clock_14_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_14_in_endofpacket_from_sa <= nios2_clock_14_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_14_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_14_in;
  --cpu_0/data_master saved-grant nios2_clock_14/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_14_in <= internal_cpu_0_data_master_requests_nios2_clock_14_in;
  --allow new arb cycle for nios2_clock_14/in, which is an e_assign
  nios2_clock_14_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_14_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_14_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_14_in_reset_n assignment, which is an e_assign
  nios2_clock_14_in_reset_n <= reset_n;
  --nios2_clock_14_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_14_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_14_in_begins_xfer) = '1'), nios2_clock_14_in_unreg_firsttransfer, nios2_clock_14_in_reg_firsttransfer);
  --nios2_clock_14_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_14_in_unreg_firsttransfer <= NOT ((nios2_clock_14_in_slavearbiterlockenable AND nios2_clock_14_in_any_continuerequest));
  --nios2_clock_14_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_14_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_14_in_begins_xfer) = '1' then 
        nios2_clock_14_in_reg_firsttransfer <= nios2_clock_14_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_14_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_14_in_beginbursttransfer_internal <= nios2_clock_14_in_begins_xfer;
  --nios2_clock_14_in_read assignment, which is an e_mux
  nios2_clock_14_in_read <= internal_cpu_0_data_master_granted_nios2_clock_14_in AND cpu_0_data_master_read;
  --nios2_clock_14_in_write assignment, which is an e_mux
  nios2_clock_14_in_write <= ((internal_cpu_0_data_master_granted_nios2_clock_14_in AND cpu_0_data_master_write)) AND nios2_clock_14_in_pretend_byte_enable;
  shifted_address_to_nios2_clock_14_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_14_in_address mux, which is an e_mux
  nios2_clock_14_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_14_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --slaveid nios2_clock_14_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_14_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_14_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_14_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_14_in_end_xfer <= nios2_clock_14_in_end_xfer;
    end if;

  end process;

  --nios2_clock_14_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_14_in_waits_for_read <= nios2_clock_14_in_in_a_read_cycle AND internal_nios2_clock_14_in_waitrequest_from_sa;
  --nios2_clock_14_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_14_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_14_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_14_in_in_a_read_cycle;
  --nios2_clock_14_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_14_in_waits_for_write <= nios2_clock_14_in_in_a_write_cycle AND internal_nios2_clock_14_in_waitrequest_from_sa;
  --nios2_clock_14_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_14_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_14_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_14_in_in_a_write_cycle;
  wait_for_nios2_clock_14_in_counter <= std_logic'('0');
  --nios2_clock_14_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios2_clock_14_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_14_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_14_in <= internal_cpu_0_data_master_granted_nios2_clock_14_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_14_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_14_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_14_in <= internal_cpu_0_data_master_requests_nios2_clock_14_in;
  --vhdl renameroo for output signals
  nios2_clock_14_in_waitrequest_from_sa <= internal_nios2_clock_14_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_14/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_14_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_switch_pio_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_14_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_14_out_granted_switch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_14_out_qualified_request_switch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_14_out_read : IN STD_LOGIC;
                 signal nios2_clock_14_out_read_data_valid_switch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_14_out_requests_switch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_14_out_write : IN STD_LOGIC;
                 signal nios2_clock_14_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal switch_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- outputs:
                 signal nios2_clock_14_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_14_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_14_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_14_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_14_out_arbitrator;


architecture europa of nios2_clock_14_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_14_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_clock_14_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_14_out_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_14_out_run :  STD_LOGIC;
                signal nios2_clock_14_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_14_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_14_out_qualified_request_switch_pio_s1 OR NOT nios2_clock_14_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_switch_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_14_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_14_out_qualified_request_switch_pio_s1 OR NOT nios2_clock_14_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_14_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_14_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_14_out_address_to_slave <= nios2_clock_14_out_address;
  --nios2_clock_14/out readdata mux, which is an e_mux
  nios2_clock_14_out_readdata <= std_logic_vector'("0000") & (switch_pio_s1_readdata_from_sa);
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_14_out_waitrequest <= NOT nios2_clock_14_out_run;
  --nios2_clock_14_out_reset_n assignment, which is an e_assign
  nios2_clock_14_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_14_out_address_to_slave <= internal_nios2_clock_14_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_14_out_waitrequest <= internal_nios2_clock_14_out_waitrequest;
--synthesis translate_off
    --nios2_clock_14_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_14_out_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_14_out_address_last_time <= nios2_clock_14_out_address;
      end if;

    end process;

    --nios2_clock_14/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_14_out_waitrequest AND ((nios2_clock_14_out_read OR nios2_clock_14_out_write));
      end if;

    end process;

    --nios2_clock_14_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_14_out_address /= nios2_clock_14_out_address_last_time))))) = '1' then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("nios2_clock_14_out_address did not heed wait!!!"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_14_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_14_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_14_out_read_last_time <= nios2_clock_14_out_read;
      end if;

    end process;

    --nios2_clock_14_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_14_out_read) /= std_logic'(nios2_clock_14_out_read_last_time)))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("nios2_clock_14_out_read did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_14_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_14_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_14_out_write_last_time <= nios2_clock_14_out_write;
      end if;

    end process;

    --nios2_clock_14_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_14_out_write) /= std_logic'(nios2_clock_14_out_write_last_time)))))) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("nios2_clock_14_out_write did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_14_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_14_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios2_clock_14_out_writedata_last_time <= nios2_clock_14_out_writedata;
      end if;

    end process;

    --nios2_clock_14_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_14_out_writedata /= nios2_clock_14_out_writedata_last_time)))) AND nios2_clock_14_out_write)) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("nios2_clock_14_out_writedata did not heed wait!!!"));
          write(output, write_line38.all);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_15_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_15_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_15_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_15_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_15_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_15_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_15_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_15_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_15_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_15_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_15_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_15_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_15_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_15_in_read : OUT STD_LOGIC;
                 signal nios2_clock_15_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_15_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_15_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_15_in_write : OUT STD_LOGIC;
                 signal nios2_clock_15_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity nios2_clock_15_in_arbitrator;


architecture europa of nios2_clock_15_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_15_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_15_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_15_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_15_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_15_in :  STD_LOGIC;
                signal internal_nios2_clock_15_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_15_in_allgrants :  STD_LOGIC;
                signal nios2_clock_15_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_15_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_15_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_15_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_15_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_15_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_15_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_15_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_15_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_15_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_15_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_15_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_15_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_15_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_15_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_15_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_15_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_15_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_15_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_15_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_15_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_15_in_end_xfer;
    end if;

  end process;

  nios2_clock_15_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_15_in);
  --assign nios2_clock_15_in_readdata_from_sa = nios2_clock_15_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_15_in_readdata_from_sa <= nios2_clock_15_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_15_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000010100000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_15_in_waitrequest_from_sa = nios2_clock_15_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_15_in_waitrequest_from_sa <= nios2_clock_15_in_waitrequest;
  --nios2_clock_15_in_arb_share_counter set values, which is an e_mux
  nios2_clock_15_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_15_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_15_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_15_in;
  --nios2_clock_15_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_15_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_15_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_15_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_15_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_15_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_15_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_15_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_15_in_allgrants all slave grants, which is an e_mux
  nios2_clock_15_in_allgrants <= nios2_clock_15_in_grant_vector;
  --nios2_clock_15_in_end_xfer assignment, which is an e_assign
  nios2_clock_15_in_end_xfer <= NOT ((nios2_clock_15_in_waits_for_read OR nios2_clock_15_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_15_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_15_in <= nios2_clock_15_in_end_xfer AND (((NOT nios2_clock_15_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_15_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_15_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_15_in AND nios2_clock_15_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_15_in AND NOT nios2_clock_15_in_non_bursting_master_requests));
  --nios2_clock_15_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_15_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_15_in_arb_counter_enable) = '1' then 
        nios2_clock_15_in_arb_share_counter <= nios2_clock_15_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_15_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_15_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_15_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_15_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_15_in AND NOT nios2_clock_15_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_15_in_slavearbiterlockenable <= or_reduce(nios2_clock_15_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_15/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_15_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_15_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_15_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_15_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_15/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_15_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_15_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_15_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_15_in <= internal_cpu_0_data_master_requests_nios2_clock_15_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_15_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_15_in <= (internal_cpu_0_data_master_granted_nios2_clock_15_in AND cpu_0_data_master_read) AND NOT nios2_clock_15_in_waits_for_read;
  --nios2_clock_15_in_writedata mux, which is an e_mux
  nios2_clock_15_in_writedata <= cpu_0_data_master_writedata (15 DOWNTO 0);
  --assign nios2_clock_15_in_endofpacket_from_sa = nios2_clock_15_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_15_in_endofpacket_from_sa <= nios2_clock_15_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_15_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_15_in;
  --cpu_0/data_master saved-grant nios2_clock_15/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_15_in <= internal_cpu_0_data_master_requests_nios2_clock_15_in;
  --allow new arb cycle for nios2_clock_15/in, which is an e_assign
  nios2_clock_15_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_15_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_15_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_15_in_reset_n assignment, which is an e_assign
  nios2_clock_15_in_reset_n <= reset_n;
  --nios2_clock_15_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_15_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_15_in_begins_xfer) = '1'), nios2_clock_15_in_unreg_firsttransfer, nios2_clock_15_in_reg_firsttransfer);
  --nios2_clock_15_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_15_in_unreg_firsttransfer <= NOT ((nios2_clock_15_in_slavearbiterlockenable AND nios2_clock_15_in_any_continuerequest));
  --nios2_clock_15_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_15_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_15_in_begins_xfer) = '1' then 
        nios2_clock_15_in_reg_firsttransfer <= nios2_clock_15_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_15_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_15_in_beginbursttransfer_internal <= nios2_clock_15_in_begins_xfer;
  --nios2_clock_15_in_read assignment, which is an e_mux
  nios2_clock_15_in_read <= internal_cpu_0_data_master_granted_nios2_clock_15_in AND cpu_0_data_master_read;
  --nios2_clock_15_in_write assignment, which is an e_mux
  nios2_clock_15_in_write <= internal_cpu_0_data_master_granted_nios2_clock_15_in AND cpu_0_data_master_write;
  shifted_address_to_nios2_clock_15_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_15_in_address mux, which is an e_mux
  nios2_clock_15_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_15_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --slaveid nios2_clock_15_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_15_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_15_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_15_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_15_in_end_xfer <= nios2_clock_15_in_end_xfer;
    end if;

  end process;

  --nios2_clock_15_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_15_in_waits_for_read <= nios2_clock_15_in_in_a_read_cycle AND internal_nios2_clock_15_in_waitrequest_from_sa;
  --nios2_clock_15_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_15_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_15_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_15_in_in_a_read_cycle;
  --nios2_clock_15_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_15_in_waits_for_write <= nios2_clock_15_in_in_a_write_cycle AND internal_nios2_clock_15_in_waitrequest_from_sa;
  --nios2_clock_15_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_15_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_15_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_15_in_in_a_write_cycle;
  wait_for_nios2_clock_15_in_counter <= std_logic'('0');
  --nios2_clock_15_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_15_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_15_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_15_in <= internal_cpu_0_data_master_granted_nios2_clock_15_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_15_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_15_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_15_in <= internal_cpu_0_data_master_requests_nios2_clock_15_in;
  --vhdl renameroo for output signals
  nios2_clock_15_in_waitrequest_from_sa <= internal_nios2_clock_15_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_15/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_15_out_arbitrator is 
        port (
              -- inputs:
                 signal cal_dac_code_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_cal_dac_code_pio_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_15_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_15_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_15_out_granted_cal_dac_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_15_out_read : IN STD_LOGIC;
                 signal nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_15_out_requests_cal_dac_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_15_out_write : IN STD_LOGIC;
                 signal nios2_clock_15_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_15_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_15_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_15_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_15_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_15_out_arbitrator;


architecture europa of nios2_clock_15_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_15_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_nios2_clock_15_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_15_out_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_15_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_15_out_run :  STD_LOGIC;
                signal nios2_clock_15_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_15_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 OR NOT nios2_clock_15_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cal_dac_code_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_15_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 OR NOT nios2_clock_15_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_15_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_15_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_15_out_address_to_slave <= nios2_clock_15_out_address;
  --nios2_clock_15/out readdata mux, which is an e_mux
  nios2_clock_15_out_readdata <= std_logic_vector'("00") & (cal_dac_code_pio_s1_readdata_from_sa);
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_15_out_waitrequest <= NOT nios2_clock_15_out_run;
  --nios2_clock_15_out_reset_n assignment, which is an e_assign
  nios2_clock_15_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_15_out_address_to_slave <= internal_nios2_clock_15_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_15_out_waitrequest <= internal_nios2_clock_15_out_waitrequest;
--synthesis translate_off
    --nios2_clock_15_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_15_out_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        nios2_clock_15_out_address_last_time <= nios2_clock_15_out_address;
      end if;

    end process;

    --nios2_clock_15/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_15_out_waitrequest AND ((nios2_clock_15_out_read OR nios2_clock_15_out_write));
      end if;

    end process;

    --nios2_clock_15_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_15_out_address /= nios2_clock_15_out_address_last_time))))) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("nios2_clock_15_out_address did not heed wait!!!"));
          write(output, write_line39.all);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_15_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_15_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_15_out_byteenable_last_time <= nios2_clock_15_out_byteenable;
      end if;

    end process;

    --nios2_clock_15_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_15_out_byteenable /= nios2_clock_15_out_byteenable_last_time))))) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("nios2_clock_15_out_byteenable did not heed wait!!!"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_15_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_15_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_15_out_read_last_time <= nios2_clock_15_out_read;
      end if;

    end process;

    --nios2_clock_15_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_15_out_read) /= std_logic'(nios2_clock_15_out_read_last_time)))))) = '1' then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("nios2_clock_15_out_read did not heed wait!!!"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_15_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_15_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_15_out_write_last_time <= nios2_clock_15_out_write;
      end if;

    end process;

    --nios2_clock_15_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_15_out_write) /= std_logic'(nios2_clock_15_out_write_last_time)))))) = '1' then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("nios2_clock_15_out_write did not heed wait!!!"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_15_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_15_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_15_out_writedata_last_time <= nios2_clock_15_out_writedata;
      end if;

    end process;

    --nios2_clock_15_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_15_out_writedata /= nios2_clock_15_out_writedata_last_time)))) AND nios2_clock_15_out_write)) = '1' then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("nios2_clock_15_out_writedata did not heed wait!!!"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_16_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_16_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_16_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_16_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_16_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_16_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_16_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_16_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_16_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_16_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_16_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_16_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_16_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_16_in_read : OUT STD_LOGIC;
                 signal nios2_clock_16_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_16_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_16_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_16_in_write : OUT STD_LOGIC;
                 signal nios2_clock_16_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_clock_16_in_arbitrator;


architecture europa of nios2_clock_16_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_16_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_16_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_16_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_16_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_16_in :  STD_LOGIC;
                signal internal_nios2_clock_16_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_16_in_allgrants :  STD_LOGIC;
                signal nios2_clock_16_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_16_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_16_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_16_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_16_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_16_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_16_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_16_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_16_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_16_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_16_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_16_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_16_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_16_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_16_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_16_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_16_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_16_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_16_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_16_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_16_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_16_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_16_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_16_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_16_in_end_xfer;
    end if;

  end process;

  nios2_clock_16_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_16_in);
  --assign nios2_clock_16_in_readdata_from_sa = nios2_clock_16_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_16_in_readdata_from_sa <= nios2_clock_16_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_16_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000010110000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_16_in_waitrequest_from_sa = nios2_clock_16_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_16_in_waitrequest_from_sa <= nios2_clock_16_in_waitrequest;
  --nios2_clock_16_in_arb_share_counter set values, which is an e_mux
  nios2_clock_16_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_16_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_16_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_16_in;
  --nios2_clock_16_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_16_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_16_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_16_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_16_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_16_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_16_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_16_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_16_in_allgrants all slave grants, which is an e_mux
  nios2_clock_16_in_allgrants <= nios2_clock_16_in_grant_vector;
  --nios2_clock_16_in_end_xfer assignment, which is an e_assign
  nios2_clock_16_in_end_xfer <= NOT ((nios2_clock_16_in_waits_for_read OR nios2_clock_16_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_16_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_16_in <= nios2_clock_16_in_end_xfer AND (((NOT nios2_clock_16_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_16_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_16_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_16_in AND nios2_clock_16_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_16_in AND NOT nios2_clock_16_in_non_bursting_master_requests));
  --nios2_clock_16_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_16_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_16_in_arb_counter_enable) = '1' then 
        nios2_clock_16_in_arb_share_counter <= nios2_clock_16_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_16_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_16_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_16_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_16_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_16_in AND NOT nios2_clock_16_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_16_in_slavearbiterlockenable <= or_reduce(nios2_clock_16_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_16/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_16_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_16_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_16_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_16_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_16/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_16_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_16_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_16_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_16_in <= internal_cpu_0_data_master_requests_nios2_clock_16_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_16_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_16_in <= (internal_cpu_0_data_master_granted_nios2_clock_16_in AND cpu_0_data_master_read) AND NOT nios2_clock_16_in_waits_for_read;
  --nios2_clock_16_in_writedata mux, which is an e_mux
  nios2_clock_16_in_writedata <= cpu_0_data_master_writedata;
  --assign nios2_clock_16_in_endofpacket_from_sa = nios2_clock_16_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_16_in_endofpacket_from_sa <= nios2_clock_16_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_16_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_16_in;
  --cpu_0/data_master saved-grant nios2_clock_16/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_16_in <= internal_cpu_0_data_master_requests_nios2_clock_16_in;
  --allow new arb cycle for nios2_clock_16/in, which is an e_assign
  nios2_clock_16_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_16_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_16_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_16_in_reset_n assignment, which is an e_assign
  nios2_clock_16_in_reset_n <= reset_n;
  --nios2_clock_16_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_16_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_16_in_begins_xfer) = '1'), nios2_clock_16_in_unreg_firsttransfer, nios2_clock_16_in_reg_firsttransfer);
  --nios2_clock_16_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_16_in_unreg_firsttransfer <= NOT ((nios2_clock_16_in_slavearbiterlockenable AND nios2_clock_16_in_any_continuerequest));
  --nios2_clock_16_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_16_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_16_in_begins_xfer) = '1' then 
        nios2_clock_16_in_reg_firsttransfer <= nios2_clock_16_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_16_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_16_in_beginbursttransfer_internal <= nios2_clock_16_in_begins_xfer;
  --nios2_clock_16_in_read assignment, which is an e_mux
  nios2_clock_16_in_read <= internal_cpu_0_data_master_granted_nios2_clock_16_in AND cpu_0_data_master_read;
  --nios2_clock_16_in_write assignment, which is an e_mux
  nios2_clock_16_in_write <= internal_cpu_0_data_master_granted_nios2_clock_16_in AND cpu_0_data_master_write;
  shifted_address_to_nios2_clock_16_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_16_in_address mux, which is an e_mux
  nios2_clock_16_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_16_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --slaveid nios2_clock_16_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_16_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_16_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_16_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_16_in_end_xfer <= nios2_clock_16_in_end_xfer;
    end if;

  end process;

  --nios2_clock_16_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_16_in_waits_for_read <= nios2_clock_16_in_in_a_read_cycle AND internal_nios2_clock_16_in_waitrequest_from_sa;
  --nios2_clock_16_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_16_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_16_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_16_in_in_a_read_cycle;
  --nios2_clock_16_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_16_in_waits_for_write <= nios2_clock_16_in_in_a_write_cycle AND internal_nios2_clock_16_in_waitrequest_from_sa;
  --nios2_clock_16_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_16_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_16_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_16_in_in_a_write_cycle;
  wait_for_nios2_clock_16_in_counter <= std_logic'('0');
  --nios2_clock_16_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_16_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_16_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_16_in <= internal_cpu_0_data_master_granted_nios2_clock_16_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_16_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_16_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_16_in <= internal_cpu_0_data_master_requests_nios2_clock_16_in;
  --vhdl renameroo for output signals
  nios2_clock_16_in_waitrequest_from_sa <= internal_nios2_clock_16_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_16/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_16_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_usb_code_pio_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_16_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_16_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_16_out_granted_usb_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_16_out_qualified_request_usb_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_16_out_read : IN STD_LOGIC;
                 signal nios2_clock_16_out_read_data_valid_usb_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_16_out_requests_usb_code_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_16_out_write : IN STD_LOGIC;
                 signal nios2_clock_16_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal usb_code_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (20 DOWNTO 0);

              -- outputs:
                 signal nios2_clock_16_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_16_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_16_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_16_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_16_out_arbitrator;


architecture europa of nios2_clock_16_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_16_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_clock_16_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_16_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_16_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_16_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_16_out_run :  STD_LOGIC;
                signal nios2_clock_16_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_16_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_16_out_qualified_request_usb_code_pio_s1 OR NOT nios2_clock_16_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_usb_code_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_16_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_16_out_qualified_request_usb_code_pio_s1 OR NOT nios2_clock_16_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_16_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_16_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_16_out_address_to_slave <= nios2_clock_16_out_address;
  --nios2_clock_16/out readdata mux, which is an e_mux
  nios2_clock_16_out_readdata <= std_logic_vector'("00000000000") & (usb_code_pio_s1_readdata_from_sa);
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_16_out_waitrequest <= NOT nios2_clock_16_out_run;
  --nios2_clock_16_out_reset_n assignment, which is an e_assign
  nios2_clock_16_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_16_out_address_to_slave <= internal_nios2_clock_16_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_16_out_waitrequest <= internal_nios2_clock_16_out_waitrequest;
--synthesis translate_off
    --nios2_clock_16_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_16_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_16_out_address_last_time <= nios2_clock_16_out_address;
      end if;

    end process;

    --nios2_clock_16/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_16_out_waitrequest AND ((nios2_clock_16_out_read OR nios2_clock_16_out_write));
      end if;

    end process;

    --nios2_clock_16_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_16_out_address /= nios2_clock_16_out_address_last_time))))) = '1' then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("nios2_clock_16_out_address did not heed wait!!!"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_16_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_16_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_16_out_byteenable_last_time <= nios2_clock_16_out_byteenable;
      end if;

    end process;

    --nios2_clock_16_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_16_out_byteenable /= nios2_clock_16_out_byteenable_last_time))))) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("nios2_clock_16_out_byteenable did not heed wait!!!"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_16_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_16_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_16_out_read_last_time <= nios2_clock_16_out_read;
      end if;

    end process;

    --nios2_clock_16_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_16_out_read) /= std_logic'(nios2_clock_16_out_read_last_time)))))) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("nios2_clock_16_out_read did not heed wait!!!"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_16_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_16_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_16_out_write_last_time <= nios2_clock_16_out_write;
      end if;

    end process;

    --nios2_clock_16_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_16_out_write) /= std_logic'(nios2_clock_16_out_write_last_time)))))) = '1' then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("nios2_clock_16_out_write did not heed wait!!!"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_16_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_16_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_16_out_writedata_last_time <= nios2_clock_16_out_writedata;
      end if;

    end process;

    --nios2_clock_16_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_16_out_writedata /= nios2_clock_16_out_writedata_last_time)))) AND nios2_clock_16_out_write)) = '1' then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("nios2_clock_16_out_writedata did not heed wait!!!"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_17_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_17_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_17_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_17_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_17_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_17_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_17_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_17_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_17_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_17_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_17_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_17_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_17_in_read : OUT STD_LOGIC;
                 signal nios2_clock_17_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_17_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_17_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_17_in_write : OUT STD_LOGIC;
                 signal nios2_clock_17_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios2_clock_17_in_arbitrator;


architecture europa of nios2_clock_17_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_17_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_17_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_17_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_17_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_17_in :  STD_LOGIC;
                signal internal_nios2_clock_17_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_17_in_allgrants :  STD_LOGIC;
                signal nios2_clock_17_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_17_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_17_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_17_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_17_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_17_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_17_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_17_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_17_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_17_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_17_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_17_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_17_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_17_in_pretend_byte_enable :  STD_LOGIC;
                signal nios2_clock_17_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_17_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_17_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_17_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_17_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_17_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_17_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_17_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_17_in_end_xfer;
    end if;

  end process;

  nios2_clock_17_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_17_in);
  --assign nios2_clock_17_in_readdata_from_sa = nios2_clock_17_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_17_in_readdata_from_sa <= nios2_clock_17_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_17_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000011000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_17_in_waitrequest_from_sa = nios2_clock_17_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_17_in_waitrequest_from_sa <= nios2_clock_17_in_waitrequest;
  --nios2_clock_17_in_arb_share_counter set values, which is an e_mux
  nios2_clock_17_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_17_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_17_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_17_in;
  --nios2_clock_17_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_17_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_17_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_17_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_17_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_17_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_17_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_17_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_17_in_allgrants all slave grants, which is an e_mux
  nios2_clock_17_in_allgrants <= nios2_clock_17_in_grant_vector;
  --nios2_clock_17_in_end_xfer assignment, which is an e_assign
  nios2_clock_17_in_end_xfer <= NOT ((nios2_clock_17_in_waits_for_read OR nios2_clock_17_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_17_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_17_in <= nios2_clock_17_in_end_xfer AND (((NOT nios2_clock_17_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_17_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_17_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_17_in AND nios2_clock_17_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_17_in AND NOT nios2_clock_17_in_non_bursting_master_requests));
  --nios2_clock_17_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_17_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_17_in_arb_counter_enable) = '1' then 
        nios2_clock_17_in_arb_share_counter <= nios2_clock_17_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_17_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_17_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_17_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_17_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_17_in AND NOT nios2_clock_17_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_17_in_slavearbiterlockenable <= or_reduce(nios2_clock_17_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_17/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_17_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_17_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_17_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_17_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_17/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_17_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_17_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_17_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_17_in <= internal_cpu_0_data_master_requests_nios2_clock_17_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_17_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_17_in <= (internal_cpu_0_data_master_granted_nios2_clock_17_in AND cpu_0_data_master_read) AND NOT nios2_clock_17_in_waits_for_read;
  --nios2_clock_17_in_writedata mux, which is an e_mux
  nios2_clock_17_in_writedata <= cpu_0_data_master_writedata (7 DOWNTO 0);
  --assign nios2_clock_17_in_endofpacket_from_sa = nios2_clock_17_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_17_in_endofpacket_from_sa <= nios2_clock_17_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_17_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_17_in;
  --cpu_0/data_master saved-grant nios2_clock_17/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_17_in <= internal_cpu_0_data_master_requests_nios2_clock_17_in;
  --allow new arb cycle for nios2_clock_17/in, which is an e_assign
  nios2_clock_17_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_17_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_17_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_17_in_reset_n assignment, which is an e_assign
  nios2_clock_17_in_reset_n <= reset_n;
  --nios2_clock_17_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_17_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_17_in_begins_xfer) = '1'), nios2_clock_17_in_unreg_firsttransfer, nios2_clock_17_in_reg_firsttransfer);
  --nios2_clock_17_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_17_in_unreg_firsttransfer <= NOT ((nios2_clock_17_in_slavearbiterlockenable AND nios2_clock_17_in_any_continuerequest));
  --nios2_clock_17_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_17_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_17_in_begins_xfer) = '1' then 
        nios2_clock_17_in_reg_firsttransfer <= nios2_clock_17_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_17_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_17_in_beginbursttransfer_internal <= nios2_clock_17_in_begins_xfer;
  --nios2_clock_17_in_read assignment, which is an e_mux
  nios2_clock_17_in_read <= internal_cpu_0_data_master_granted_nios2_clock_17_in AND cpu_0_data_master_read;
  --nios2_clock_17_in_write assignment, which is an e_mux
  nios2_clock_17_in_write <= ((internal_cpu_0_data_master_granted_nios2_clock_17_in AND cpu_0_data_master_write)) AND nios2_clock_17_in_pretend_byte_enable;
  shifted_address_to_nios2_clock_17_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_17_in_address mux, which is an e_mux
  nios2_clock_17_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_17_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --slaveid nios2_clock_17_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_17_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_17_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_17_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_17_in_end_xfer <= nios2_clock_17_in_end_xfer;
    end if;

  end process;

  --nios2_clock_17_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_17_in_waits_for_read <= nios2_clock_17_in_in_a_read_cycle AND internal_nios2_clock_17_in_waitrequest_from_sa;
  --nios2_clock_17_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_17_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_17_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_17_in_in_a_read_cycle;
  --nios2_clock_17_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_17_in_waits_for_write <= nios2_clock_17_in_in_a_write_cycle AND internal_nios2_clock_17_in_waitrequest_from_sa;
  --nios2_clock_17_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_17_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_17_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_17_in_in_a_write_cycle;
  wait_for_nios2_clock_17_in_counter <= std_logic'('0');
  --nios2_clock_17_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios2_clock_17_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_17_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_17_in <= internal_cpu_0_data_master_granted_nios2_clock_17_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_17_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_17_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_17_in <= internal_cpu_0_data_master_requests_nios2_clock_17_in;
  --vhdl renameroo for output signals
  nios2_clock_17_in_waitrequest_from_sa <= internal_nios2_clock_17_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_17/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_17_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sample_and_hold_pio_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_17_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_17_out_granted_sample_and_hold_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_17_out_read : IN STD_LOGIC;
                 signal nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_17_out_requests_sample_and_hold_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_17_out_write : IN STD_LOGIC;
                 signal nios2_clock_17_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sample_and_hold_pio_s1_readdata_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_17_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_17_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_17_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_17_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_17_out_arbitrator;


architecture europa of nios2_clock_17_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_17_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_clock_17_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_17_out_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_17_out_run :  STD_LOGIC;
                signal nios2_clock_17_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_17_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 OR NOT nios2_clock_17_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sample_and_hold_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_17_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 OR NOT nios2_clock_17_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_17_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_17_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_17_out_address_to_slave <= nios2_clock_17_out_address;
  --nios2_clock_17/out readdata mux, which is an e_mux
  nios2_clock_17_out_readdata <= std_logic_vector'("0000000") & (A_TOSTDLOGICVECTOR(sample_and_hold_pio_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_17_out_waitrequest <= NOT nios2_clock_17_out_run;
  --nios2_clock_17_out_reset_n assignment, which is an e_assign
  nios2_clock_17_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_17_out_address_to_slave <= internal_nios2_clock_17_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_17_out_waitrequest <= internal_nios2_clock_17_out_waitrequest;
--synthesis translate_off
    --nios2_clock_17_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_17_out_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_17_out_address_last_time <= nios2_clock_17_out_address;
      end if;

    end process;

    --nios2_clock_17/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_17_out_waitrequest AND ((nios2_clock_17_out_read OR nios2_clock_17_out_write));
      end if;

    end process;

    --nios2_clock_17_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_17_out_address /= nios2_clock_17_out_address_last_time))))) = '1' then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("nios2_clock_17_out_address did not heed wait!!!"));
          write(output, write_line49.all);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_17_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_17_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_17_out_read_last_time <= nios2_clock_17_out_read;
      end if;

    end process;

    --nios2_clock_17_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_17_out_read) /= std_logic'(nios2_clock_17_out_read_last_time)))))) = '1' then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("nios2_clock_17_out_read did not heed wait!!!"));
          write(output, write_line50.all);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_17_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_17_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_17_out_write_last_time <= nios2_clock_17_out_write;
      end if;

    end process;

    --nios2_clock_17_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_17_out_write) /= std_logic'(nios2_clock_17_out_write_last_time)))))) = '1' then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("nios2_clock_17_out_write did not heed wait!!!"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_17_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_17_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios2_clock_17_out_writedata_last_time <= nios2_clock_17_out_writedata;
      end if;

    end process;

    --nios2_clock_17_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_17_out_writedata /= nios2_clock_17_out_writedata_last_time)))) AND nios2_clock_17_out_write)) = '1' then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("nios2_clock_17_out_writedata did not heed wait!!!"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_18_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_18_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_18_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_18_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_18_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_18_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_18_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_18_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_18_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_18_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_18_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_18_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_18_in_read : OUT STD_LOGIC;
                 signal nios2_clock_18_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_18_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_18_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_18_in_write : OUT STD_LOGIC;
                 signal nios2_clock_18_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity nios2_clock_18_in_arbitrator;


architecture europa of nios2_clock_18_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_18_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_18_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_18_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_18_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_18_in :  STD_LOGIC;
                signal internal_nios2_clock_18_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_18_in_allgrants :  STD_LOGIC;
                signal nios2_clock_18_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_18_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_18_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_18_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_18_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_18_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_18_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_18_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_18_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_18_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_18_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_18_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_18_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_18_in_pretend_byte_enable :  STD_LOGIC;
                signal nios2_clock_18_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_18_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_18_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_18_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_18_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_18_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_18_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_18_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_18_in_end_xfer;
    end if;

  end process;

  nios2_clock_18_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_18_in);
  --assign nios2_clock_18_in_readdata_from_sa = nios2_clock_18_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_18_in_readdata_from_sa <= nios2_clock_18_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_18_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000011010000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_18_in_waitrequest_from_sa = nios2_clock_18_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_18_in_waitrequest_from_sa <= nios2_clock_18_in_waitrequest;
  --nios2_clock_18_in_arb_share_counter set values, which is an e_mux
  nios2_clock_18_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_18_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_18_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_18_in;
  --nios2_clock_18_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_18_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_18_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_18_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_18_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_18_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_18_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_18_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_18_in_allgrants all slave grants, which is an e_mux
  nios2_clock_18_in_allgrants <= nios2_clock_18_in_grant_vector;
  --nios2_clock_18_in_end_xfer assignment, which is an e_assign
  nios2_clock_18_in_end_xfer <= NOT ((nios2_clock_18_in_waits_for_read OR nios2_clock_18_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_18_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_18_in <= nios2_clock_18_in_end_xfer AND (((NOT nios2_clock_18_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_18_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_18_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_18_in AND nios2_clock_18_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_18_in AND NOT nios2_clock_18_in_non_bursting_master_requests));
  --nios2_clock_18_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_18_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_18_in_arb_counter_enable) = '1' then 
        nios2_clock_18_in_arb_share_counter <= nios2_clock_18_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_18_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_18_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_18_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_18_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_18_in AND NOT nios2_clock_18_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_18_in_slavearbiterlockenable <= or_reduce(nios2_clock_18_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_18/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_18_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_18_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_18_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_18_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_18/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_18_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_18_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_18_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_18_in <= internal_cpu_0_data_master_requests_nios2_clock_18_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_18_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_18_in <= (internal_cpu_0_data_master_granted_nios2_clock_18_in AND cpu_0_data_master_read) AND NOT nios2_clock_18_in_waits_for_read;
  --nios2_clock_18_in_writedata mux, which is an e_mux
  nios2_clock_18_in_writedata <= cpu_0_data_master_writedata (7 DOWNTO 0);
  --assign nios2_clock_18_in_endofpacket_from_sa = nios2_clock_18_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_18_in_endofpacket_from_sa <= nios2_clock_18_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_18_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_18_in;
  --cpu_0/data_master saved-grant nios2_clock_18/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_18_in <= internal_cpu_0_data_master_requests_nios2_clock_18_in;
  --allow new arb cycle for nios2_clock_18/in, which is an e_assign
  nios2_clock_18_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_18_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_18_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_18_in_reset_n assignment, which is an e_assign
  nios2_clock_18_in_reset_n <= reset_n;
  --nios2_clock_18_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_18_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_18_in_begins_xfer) = '1'), nios2_clock_18_in_unreg_firsttransfer, nios2_clock_18_in_reg_firsttransfer);
  --nios2_clock_18_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_18_in_unreg_firsttransfer <= NOT ((nios2_clock_18_in_slavearbiterlockenable AND nios2_clock_18_in_any_continuerequest));
  --nios2_clock_18_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_18_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_18_in_begins_xfer) = '1' then 
        nios2_clock_18_in_reg_firsttransfer <= nios2_clock_18_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_18_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_18_in_beginbursttransfer_internal <= nios2_clock_18_in_begins_xfer;
  --nios2_clock_18_in_read assignment, which is an e_mux
  nios2_clock_18_in_read <= internal_cpu_0_data_master_granted_nios2_clock_18_in AND cpu_0_data_master_read;
  --nios2_clock_18_in_write assignment, which is an e_mux
  nios2_clock_18_in_write <= ((internal_cpu_0_data_master_granted_nios2_clock_18_in AND cpu_0_data_master_write)) AND nios2_clock_18_in_pretend_byte_enable;
  shifted_address_to_nios2_clock_18_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_18_in_address mux, which is an e_mux
  nios2_clock_18_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_18_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --slaveid nios2_clock_18_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_18_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_18_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_18_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_18_in_end_xfer <= nios2_clock_18_in_end_xfer;
    end if;

  end process;

  --nios2_clock_18_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_18_in_waits_for_read <= nios2_clock_18_in_in_a_read_cycle AND internal_nios2_clock_18_in_waitrequest_from_sa;
  --nios2_clock_18_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_18_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_18_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_18_in_in_a_read_cycle;
  --nios2_clock_18_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_18_in_waits_for_write <= nios2_clock_18_in_in_a_write_cycle AND internal_nios2_clock_18_in_waitrequest_from_sa;
  --nios2_clock_18_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_18_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_18_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_18_in_in_a_write_cycle;
  wait_for_nios2_clock_18_in_counter <= std_logic'('0');
  --nios2_clock_18_in_pretend_byte_enable byte enable port mux, which is an e_mux
  nios2_clock_18_in_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_18_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_18_in <= internal_cpu_0_data_master_granted_nios2_clock_18_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_18_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_18_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_18_in <= internal_cpu_0_data_master_requests_nios2_clock_18_in;
  --vhdl renameroo for output signals
  nios2_clock_18_in_waitrequest_from_sa <= internal_nios2_clock_18_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_18/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_18_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_latch_pio_s1_end_xfer : IN STD_LOGIC;
                 signal latch_pio_s1_readdata_from_sa : IN STD_LOGIC;
                 signal nios2_clock_18_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_18_out_granted_latch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_18_out_qualified_request_latch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_18_out_read : IN STD_LOGIC;
                 signal nios2_clock_18_out_read_data_valid_latch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_18_out_requests_latch_pio_s1 : IN STD_LOGIC;
                 signal nios2_clock_18_out_write : IN STD_LOGIC;
                 signal nios2_clock_18_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_18_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_18_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_clock_18_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_18_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_18_out_arbitrator;


architecture europa of nios2_clock_18_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_18_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_clock_18_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_18_out_address_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_18_out_run :  STD_LOGIC;
                signal nios2_clock_18_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_18_out_writedata_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_18_out_qualified_request_latch_pio_s1 OR NOT nios2_clock_18_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_latch_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_18_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_18_out_qualified_request_latch_pio_s1 OR NOT nios2_clock_18_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_18_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_18_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_18_out_address_to_slave <= nios2_clock_18_out_address;
  --nios2_clock_18/out readdata mux, which is an e_mux
  nios2_clock_18_out_readdata <= std_logic_vector'("0000000") & (A_TOSTDLOGICVECTOR(latch_pio_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_18_out_waitrequest <= NOT nios2_clock_18_out_run;
  --nios2_clock_18_out_reset_n assignment, which is an e_assign
  nios2_clock_18_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_18_out_address_to_slave <= internal_nios2_clock_18_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_18_out_waitrequest <= internal_nios2_clock_18_out_waitrequest;
--synthesis translate_off
    --nios2_clock_18_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_18_out_address_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_18_out_address_last_time <= nios2_clock_18_out_address;
      end if;

    end process;

    --nios2_clock_18/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_18_out_waitrequest AND ((nios2_clock_18_out_read OR nios2_clock_18_out_write));
      end if;

    end process;

    --nios2_clock_18_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line53 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_18_out_address /= nios2_clock_18_out_address_last_time))))) = '1' then 
          write(write_line53, now);
          write(write_line53, string'(": "));
          write(write_line53, string'("nios2_clock_18_out_address did not heed wait!!!"));
          write(output, write_line53.all);
          deallocate (write_line53);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_18_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_18_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_18_out_read_last_time <= nios2_clock_18_out_read;
      end if;

    end process;

    --nios2_clock_18_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line54 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_18_out_read) /= std_logic'(nios2_clock_18_out_read_last_time)))))) = '1' then 
          write(write_line54, now);
          write(write_line54, string'(": "));
          write(write_line54, string'("nios2_clock_18_out_read did not heed wait!!!"));
          write(output, write_line54.all);
          deallocate (write_line54);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_18_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_18_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_18_out_write_last_time <= nios2_clock_18_out_write;
      end if;

    end process;

    --nios2_clock_18_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line55 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_18_out_write) /= std_logic'(nios2_clock_18_out_write_last_time)))))) = '1' then 
          write(write_line55, now);
          write(write_line55, string'(": "));
          write(write_line55, string'("nios2_clock_18_out_write did not heed wait!!!"));
          write(output, write_line55.all);
          deallocate (write_line55);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_18_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_18_out_writedata_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        nios2_clock_18_out_writedata_last_time <= nios2_clock_18_out_writedata;
      end if;

    end process;

    --nios2_clock_18_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line56 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_18_out_writedata /= nios2_clock_18_out_writedata_last_time)))) AND nios2_clock_18_out_write)) = '1' then 
          write(write_line56, now);
          write(write_line56, string'(": "));
          write(write_line56, string'("nios2_clock_18_out_writedata did not heed wait!!!"));
          write(output, write_line56.all);
          deallocate (write_line56);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_2_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_2_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_2_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_2_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_2_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_2_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_2_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_2_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_2_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_2_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_2_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_2_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_2_in_nativeaddress : OUT STD_LOGIC;
                 signal nios2_clock_2_in_read : OUT STD_LOGIC;
                 signal nios2_clock_2_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_2_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_2_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_2_in_write : OUT STD_LOGIC;
                 signal nios2_clock_2_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_clock_2_in_arbitrator;


architecture europa of nios2_clock_2_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_2_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_2_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_2_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_2_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_2_in :  STD_LOGIC;
                signal internal_nios2_clock_2_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_2_in_allgrants :  STD_LOGIC;
                signal nios2_clock_2_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_2_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_2_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_2_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_2_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_2_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_2_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_2_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_2_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_2_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_2_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_2_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_2_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_2_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_2_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_2_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_2_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_2_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_2_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_2_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_2_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_2_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_2_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_2_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_2_in_end_xfer;
    end if;

  end process;

  nios2_clock_2_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_2_in);
  --assign nios2_clock_2_in_readdata_from_sa = nios2_clock_2_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_2_in_readdata_from_sa <= nios2_clock_2_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_2_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("1000000010001000011100000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_2_in_waitrequest_from_sa = nios2_clock_2_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_2_in_waitrequest_from_sa <= nios2_clock_2_in_waitrequest;
  --nios2_clock_2_in_arb_share_counter set values, which is an e_mux
  nios2_clock_2_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_2_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_2_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_2_in;
  --nios2_clock_2_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_2_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_2_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_2_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_2_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_2_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_2_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_2_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_2_in_allgrants all slave grants, which is an e_mux
  nios2_clock_2_in_allgrants <= nios2_clock_2_in_grant_vector;
  --nios2_clock_2_in_end_xfer assignment, which is an e_assign
  nios2_clock_2_in_end_xfer <= NOT ((nios2_clock_2_in_waits_for_read OR nios2_clock_2_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_2_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_2_in <= nios2_clock_2_in_end_xfer AND (((NOT nios2_clock_2_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_2_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_2_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_2_in AND nios2_clock_2_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_2_in AND NOT nios2_clock_2_in_non_bursting_master_requests));
  --nios2_clock_2_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_2_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_2_in_arb_counter_enable) = '1' then 
        nios2_clock_2_in_arb_share_counter <= nios2_clock_2_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_2_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_2_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_2_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_2_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_2_in AND NOT nios2_clock_2_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_2_in_slavearbiterlockenable <= or_reduce(nios2_clock_2_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_2/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_2_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_2_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_2_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_2_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_2/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_2_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_2_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_2_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_2_in <= internal_cpu_0_data_master_requests_nios2_clock_2_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_2_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_2_in <= (internal_cpu_0_data_master_granted_nios2_clock_2_in AND cpu_0_data_master_read) AND NOT nios2_clock_2_in_waits_for_read;
  --nios2_clock_2_in_writedata mux, which is an e_mux
  nios2_clock_2_in_writedata <= cpu_0_data_master_writedata;
  --assign nios2_clock_2_in_endofpacket_from_sa = nios2_clock_2_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_2_in_endofpacket_from_sa <= nios2_clock_2_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_2_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_2_in;
  --cpu_0/data_master saved-grant nios2_clock_2/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_2_in <= internal_cpu_0_data_master_requests_nios2_clock_2_in;
  --allow new arb cycle for nios2_clock_2/in, which is an e_assign
  nios2_clock_2_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_2_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_2_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_2_in_reset_n assignment, which is an e_assign
  nios2_clock_2_in_reset_n <= reset_n;
  --nios2_clock_2_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_2_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_2_in_begins_xfer) = '1'), nios2_clock_2_in_unreg_firsttransfer, nios2_clock_2_in_reg_firsttransfer);
  --nios2_clock_2_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_2_in_unreg_firsttransfer <= NOT ((nios2_clock_2_in_slavearbiterlockenable AND nios2_clock_2_in_any_continuerequest));
  --nios2_clock_2_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_2_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_2_in_begins_xfer) = '1' then 
        nios2_clock_2_in_reg_firsttransfer <= nios2_clock_2_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_2_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_2_in_beginbursttransfer_internal <= nios2_clock_2_in_begins_xfer;
  --nios2_clock_2_in_read assignment, which is an e_mux
  nios2_clock_2_in_read <= internal_cpu_0_data_master_granted_nios2_clock_2_in AND cpu_0_data_master_read;
  --nios2_clock_2_in_write assignment, which is an e_mux
  nios2_clock_2_in_write <= internal_cpu_0_data_master_granted_nios2_clock_2_in AND cpu_0_data_master_write;
  shifted_address_to_nios2_clock_2_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_2_in_address mux, which is an e_mux
  nios2_clock_2_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_2_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --slaveid nios2_clock_2_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_2_in_nativeaddress <= Vector_To_Std_Logic(A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")));
  --d1_nios2_clock_2_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_2_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_2_in_end_xfer <= nios2_clock_2_in_end_xfer;
    end if;

  end process;

  --nios2_clock_2_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_2_in_waits_for_read <= nios2_clock_2_in_in_a_read_cycle AND internal_nios2_clock_2_in_waitrequest_from_sa;
  --nios2_clock_2_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_2_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_2_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_2_in_in_a_read_cycle;
  --nios2_clock_2_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_2_in_waits_for_write <= nios2_clock_2_in_in_a_write_cycle AND internal_nios2_clock_2_in_waitrequest_from_sa;
  --nios2_clock_2_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_2_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_2_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_2_in_in_a_write_cycle;
  wait_for_nios2_clock_2_in_counter <= std_logic'('0');
  --nios2_clock_2_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_2_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_2_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_2_in <= internal_cpu_0_data_master_granted_nios2_clock_2_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_2_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_2_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_2_in <= internal_cpu_0_data_master_requests_nios2_clock_2_in;
  --vhdl renameroo for output signals
  nios2_clock_2_in_waitrequest_from_sa <= internal_nios2_clock_2_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_2/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_2_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_clock_2_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal nios2_clock_2_out_read : IN STD_LOGIC;
                 signal nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal nios2_clock_2_out_write : IN STD_LOGIC;
                 signal nios2_clock_2_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_2_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_2_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_2_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_2_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_2_out_arbitrator;


architecture europa of nios2_clock_2_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_2_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_nios2_clock_2_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_2_out_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_2_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_2_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_2_out_run :  STD_LOGIC;
                signal nios2_clock_2_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_2_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave OR NOT ((nios2_clock_2_out_read OR nios2_clock_2_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_2_out_read OR nios2_clock_2_out_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave OR NOT ((nios2_clock_2_out_read OR nios2_clock_2_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_2_out_read OR nios2_clock_2_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_2_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_2_out_address_to_slave <= nios2_clock_2_out_address;
  --nios2_clock_2/out readdata mux, which is an e_mux
  nios2_clock_2_out_readdata <= jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_2_out_waitrequest <= NOT nios2_clock_2_out_run;
  --nios2_clock_2_out_reset_n assignment, which is an e_assign
  nios2_clock_2_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_2_out_address_to_slave <= internal_nios2_clock_2_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_2_out_waitrequest <= internal_nios2_clock_2_out_waitrequest;
--synthesis translate_off
    --nios2_clock_2_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_2_out_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        nios2_clock_2_out_address_last_time <= nios2_clock_2_out_address;
      end if;

    end process;

    --nios2_clock_2/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_2_out_waitrequest AND ((nios2_clock_2_out_read OR nios2_clock_2_out_write));
      end if;

    end process;

    --nios2_clock_2_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line57 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_2_out_address /= nios2_clock_2_out_address_last_time))))) = '1' then 
          write(write_line57, now);
          write(write_line57, string'(": "));
          write(write_line57, string'("nios2_clock_2_out_address did not heed wait!!!"));
          write(output, write_line57.all);
          deallocate (write_line57);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_2_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_2_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_2_out_byteenable_last_time <= nios2_clock_2_out_byteenable;
      end if;

    end process;

    --nios2_clock_2_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line58 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_2_out_byteenable /= nios2_clock_2_out_byteenable_last_time))))) = '1' then 
          write(write_line58, now);
          write(write_line58, string'(": "));
          write(write_line58, string'("nios2_clock_2_out_byteenable did not heed wait!!!"));
          write(output, write_line58.all);
          deallocate (write_line58);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_2_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_2_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_2_out_read_last_time <= nios2_clock_2_out_read;
      end if;

    end process;

    --nios2_clock_2_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line59 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_2_out_read) /= std_logic'(nios2_clock_2_out_read_last_time)))))) = '1' then 
          write(write_line59, now);
          write(write_line59, string'(": "));
          write(write_line59, string'("nios2_clock_2_out_read did not heed wait!!!"));
          write(output, write_line59.all);
          deallocate (write_line59);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_2_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_2_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_2_out_write_last_time <= nios2_clock_2_out_write;
      end if;

    end process;

    --nios2_clock_2_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line60 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_2_out_write) /= std_logic'(nios2_clock_2_out_write_last_time)))))) = '1' then 
          write(write_line60, now);
          write(write_line60, string'(": "));
          write(write_line60, string'("nios2_clock_2_out_write did not heed wait!!!"));
          write(output, write_line60.all);
          deallocate (write_line60);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_2_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_2_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_2_out_writedata_last_time <= nios2_clock_2_out_writedata;
      end if;

    end process;

    --nios2_clock_2_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line61 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_2_out_writedata /= nios2_clock_2_out_writedata_last_time)))) AND nios2_clock_2_out_write)) = '1' then 
          write(write_line61, now);
          write(write_line61, string'(": "));
          write(write_line61, string'("nios2_clock_2_out_writedata did not heed wait!!!"));
          write(output, write_line61.all);
          deallocate (write_line61);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_3_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_3_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_3_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_3_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_3_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_3_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_3_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_3_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_3_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_3_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_3_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_3_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_3_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_3_in_read : OUT STD_LOGIC;
                 signal nios2_clock_3_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_3_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_3_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_3_in_write : OUT STD_LOGIC;
                 signal nios2_clock_3_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity nios2_clock_3_in_arbitrator;


architecture europa of nios2_clock_3_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_3_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_3_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_3_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_3_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_3_in :  STD_LOGIC;
                signal internal_nios2_clock_3_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_3_in_allgrants :  STD_LOGIC;
                signal nios2_clock_3_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_3_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_3_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_3_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_3_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_3_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_3_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_3_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_3_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_3_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_3_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_3_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_3_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_3_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_3_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_3_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_3_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_3_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_3_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_3_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_3_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_3_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_3_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_3_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_3_in_end_xfer;
    end if;

  end process;

  nios2_clock_3_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_3_in);
  --assign nios2_clock_3_in_readdata_from_sa = nios2_clock_3_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_3_in_readdata_from_sa <= nios2_clock_3_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_3_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1000000010001000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_3_in_waitrequest_from_sa = nios2_clock_3_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_3_in_waitrequest_from_sa <= nios2_clock_3_in_waitrequest;
  --nios2_clock_3_in_arb_share_counter set values, which is an e_mux
  nios2_clock_3_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_3_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_3_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_3_in;
  --nios2_clock_3_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_3_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_3_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_3_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_3_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_3_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_3_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_3_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_3_in_allgrants all slave grants, which is an e_mux
  nios2_clock_3_in_allgrants <= nios2_clock_3_in_grant_vector;
  --nios2_clock_3_in_end_xfer assignment, which is an e_assign
  nios2_clock_3_in_end_xfer <= NOT ((nios2_clock_3_in_waits_for_read OR nios2_clock_3_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_3_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_3_in <= nios2_clock_3_in_end_xfer AND (((NOT nios2_clock_3_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_3_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_3_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_3_in AND nios2_clock_3_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_3_in AND NOT nios2_clock_3_in_non_bursting_master_requests));
  --nios2_clock_3_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_3_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_3_in_arb_counter_enable) = '1' then 
        nios2_clock_3_in_arb_share_counter <= nios2_clock_3_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_3_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_3_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_3_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_3_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_3_in AND NOT nios2_clock_3_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_3_in_slavearbiterlockenable <= or_reduce(nios2_clock_3_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_3/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_3_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_3_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_3_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_3_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_3/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_3_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_3_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_3_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_3_in <= internal_cpu_0_data_master_requests_nios2_clock_3_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_3_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_3_in <= (internal_cpu_0_data_master_granted_nios2_clock_3_in AND cpu_0_data_master_read) AND NOT nios2_clock_3_in_waits_for_read;
  --nios2_clock_3_in_writedata mux, which is an e_mux
  nios2_clock_3_in_writedata <= cpu_0_data_master_writedata (15 DOWNTO 0);
  --assign nios2_clock_3_in_endofpacket_from_sa = nios2_clock_3_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_3_in_endofpacket_from_sa <= nios2_clock_3_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_3_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_3_in;
  --cpu_0/data_master saved-grant nios2_clock_3/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_3_in <= internal_cpu_0_data_master_requests_nios2_clock_3_in;
  --allow new arb cycle for nios2_clock_3/in, which is an e_assign
  nios2_clock_3_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_3_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_3_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_3_in_reset_n assignment, which is an e_assign
  nios2_clock_3_in_reset_n <= reset_n;
  --nios2_clock_3_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_3_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_3_in_begins_xfer) = '1'), nios2_clock_3_in_unreg_firsttransfer, nios2_clock_3_in_reg_firsttransfer);
  --nios2_clock_3_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_3_in_unreg_firsttransfer <= NOT ((nios2_clock_3_in_slavearbiterlockenable AND nios2_clock_3_in_any_continuerequest));
  --nios2_clock_3_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_3_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_3_in_begins_xfer) = '1' then 
        nios2_clock_3_in_reg_firsttransfer <= nios2_clock_3_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_3_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_3_in_beginbursttransfer_internal <= nios2_clock_3_in_begins_xfer;
  --nios2_clock_3_in_read assignment, which is an e_mux
  nios2_clock_3_in_read <= internal_cpu_0_data_master_granted_nios2_clock_3_in AND cpu_0_data_master_read;
  --nios2_clock_3_in_write assignment, which is an e_mux
  nios2_clock_3_in_write <= internal_cpu_0_data_master_granted_nios2_clock_3_in AND cpu_0_data_master_write;
  shifted_address_to_nios2_clock_3_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_3_in_address mux, which is an e_mux
  nios2_clock_3_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_3_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --slaveid nios2_clock_3_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_3_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_nios2_clock_3_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_3_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_3_in_end_xfer <= nios2_clock_3_in_end_xfer;
    end if;

  end process;

  --nios2_clock_3_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_3_in_waits_for_read <= nios2_clock_3_in_in_a_read_cycle AND internal_nios2_clock_3_in_waitrequest_from_sa;
  --nios2_clock_3_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_3_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_3_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_3_in_in_a_read_cycle;
  --nios2_clock_3_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_3_in_waits_for_write <= nios2_clock_3_in_in_a_write_cycle AND internal_nios2_clock_3_in_waitrequest_from_sa;
  --nios2_clock_3_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_3_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_3_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_3_in_in_a_write_cycle;
  wait_for_nios2_clock_3_in_counter <= std_logic'('0');
  --nios2_clock_3_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_3_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_3_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_3_in <= internal_cpu_0_data_master_granted_nios2_clock_3_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_3_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_3_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_3_in <= internal_cpu_0_data_master_requests_nios2_clock_3_in;
  --vhdl renameroo for output signals
  nios2_clock_3_in_waitrequest_from_sa <= internal_nios2_clock_3_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_3/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_3_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_3_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_3_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_3_out_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal nios2_clock_3_out_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal nios2_clock_3_out_read : IN STD_LOGIC;
                 signal nios2_clock_3_out_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal nios2_clock_3_out_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal nios2_clock_3_out_write : IN STD_LOGIC;
                 signal nios2_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal nios2_clock_3_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_3_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_3_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_3_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_3_out_arbitrator;


architecture europa of nios2_clock_3_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_3_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_clock_3_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_3_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_3_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_3_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_3_out_run :  STD_LOGIC;
                signal nios2_clock_3_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_3_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_3_out_qualified_request_sys_clk_timer_s1 OR NOT nios2_clock_3_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sys_clk_timer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_3_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_3_out_qualified_request_sys_clk_timer_s1 OR NOT nios2_clock_3_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_3_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_3_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_3_out_address_to_slave <= nios2_clock_3_out_address;
  --nios2_clock_3/out readdata mux, which is an e_mux
  nios2_clock_3_out_readdata <= sys_clk_timer_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_3_out_waitrequest <= NOT nios2_clock_3_out_run;
  --nios2_clock_3_out_reset_n assignment, which is an e_assign
  nios2_clock_3_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_3_out_address_to_slave <= internal_nios2_clock_3_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_3_out_waitrequest <= internal_nios2_clock_3_out_waitrequest;
--synthesis translate_off
    --nios2_clock_3_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_3_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_3_out_address_last_time <= nios2_clock_3_out_address;
      end if;

    end process;

    --nios2_clock_3/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_3_out_waitrequest AND ((nios2_clock_3_out_read OR nios2_clock_3_out_write));
      end if;

    end process;

    --nios2_clock_3_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line62 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_3_out_address /= nios2_clock_3_out_address_last_time))))) = '1' then 
          write(write_line62, now);
          write(write_line62, string'(": "));
          write(write_line62, string'("nios2_clock_3_out_address did not heed wait!!!"));
          write(output, write_line62.all);
          deallocate (write_line62);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_3_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_3_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_3_out_byteenable_last_time <= nios2_clock_3_out_byteenable;
      end if;

    end process;

    --nios2_clock_3_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line63 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_3_out_byteenable /= nios2_clock_3_out_byteenable_last_time))))) = '1' then 
          write(write_line63, now);
          write(write_line63, string'(": "));
          write(write_line63, string'("nios2_clock_3_out_byteenable did not heed wait!!!"));
          write(output, write_line63.all);
          deallocate (write_line63);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_3_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_3_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_3_out_read_last_time <= nios2_clock_3_out_read;
      end if;

    end process;

    --nios2_clock_3_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line64 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_3_out_read) /= std_logic'(nios2_clock_3_out_read_last_time)))))) = '1' then 
          write(write_line64, now);
          write(write_line64, string'(": "));
          write(write_line64, string'("nios2_clock_3_out_read did not heed wait!!!"));
          write(output, write_line64.all);
          deallocate (write_line64);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_3_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_3_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_3_out_write_last_time <= nios2_clock_3_out_write;
      end if;

    end process;

    --nios2_clock_3_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line65 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_3_out_write) /= std_logic'(nios2_clock_3_out_write_last_time)))))) = '1' then 
          write(write_line65, now);
          write(write_line65, string'(": "));
          write(write_line65, string'("nios2_clock_3_out_write did not heed wait!!!"));
          write(output, write_line65.all);
          deallocate (write_line65);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_3_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_3_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_3_out_writedata_last_time <= nios2_clock_3_out_writedata;
      end if;

    end process;

    --nios2_clock_3_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line66 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_3_out_writedata /= nios2_clock_3_out_writedata_last_time)))) AND nios2_clock_3_out_write)) = '1' then 
          write(write_line66, now);
          write(write_line66, string'(": "));
          write(write_line66, string'("nios2_clock_3_out_writedata did not heed wait!!!"));
          write(output, write_line66.all);
          deallocate (write_line66);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_4_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_4_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_4_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_4_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_4_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_4_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_4_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_4_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_4_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_4_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_4_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_4_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_4_in_nativeaddress : OUT STD_LOGIC;
                 signal nios2_clock_4_in_read : OUT STD_LOGIC;
                 signal nios2_clock_4_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_4_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_4_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_4_in_write : OUT STD_LOGIC;
                 signal nios2_clock_4_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_clock_4_in_arbitrator;


architecture europa of nios2_clock_4_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_4_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_4_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_4_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_4_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_4_in :  STD_LOGIC;
                signal internal_nios2_clock_4_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_4_in_allgrants :  STD_LOGIC;
                signal nios2_clock_4_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_4_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_4_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_4_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_4_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_4_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_4_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_4_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_4_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_4_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_4_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_4_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_4_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_4_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_4_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_4_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_4_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_4_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_4_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_4_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_4_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_4_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_4_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_4_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_4_in_end_xfer;
    end if;

  end process;

  nios2_clock_4_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_4_in);
  --assign nios2_clock_4_in_readdata_from_sa = nios2_clock_4_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_4_in_readdata_from_sa <= nios2_clock_4_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_4_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("1000000010001000011101000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_4_in_waitrequest_from_sa = nios2_clock_4_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_4_in_waitrequest_from_sa <= nios2_clock_4_in_waitrequest;
  --nios2_clock_4_in_arb_share_counter set values, which is an e_mux
  nios2_clock_4_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_4_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_4_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_4_in;
  --nios2_clock_4_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_4_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_4_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_4_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_4_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_4_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_4_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_4_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_4_in_allgrants all slave grants, which is an e_mux
  nios2_clock_4_in_allgrants <= nios2_clock_4_in_grant_vector;
  --nios2_clock_4_in_end_xfer assignment, which is an e_assign
  nios2_clock_4_in_end_xfer <= NOT ((nios2_clock_4_in_waits_for_read OR nios2_clock_4_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_4_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_4_in <= nios2_clock_4_in_end_xfer AND (((NOT nios2_clock_4_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_4_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_4_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_4_in AND nios2_clock_4_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_4_in AND NOT nios2_clock_4_in_non_bursting_master_requests));
  --nios2_clock_4_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_4_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_4_in_arb_counter_enable) = '1' then 
        nios2_clock_4_in_arb_share_counter <= nios2_clock_4_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_4_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_4_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_4_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_4_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_4_in AND NOT nios2_clock_4_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_4_in_slavearbiterlockenable <= or_reduce(nios2_clock_4_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_4/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_4_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_4_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_4_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_4_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_4/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_4_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_4_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_4_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_4_in <= internal_cpu_0_data_master_requests_nios2_clock_4_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_4_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_4_in <= (internal_cpu_0_data_master_granted_nios2_clock_4_in AND cpu_0_data_master_read) AND NOT nios2_clock_4_in_waits_for_read;
  --nios2_clock_4_in_writedata mux, which is an e_mux
  nios2_clock_4_in_writedata <= cpu_0_data_master_writedata;
  --assign nios2_clock_4_in_endofpacket_from_sa = nios2_clock_4_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_4_in_endofpacket_from_sa <= nios2_clock_4_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_4_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_4_in;
  --cpu_0/data_master saved-grant nios2_clock_4/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_4_in <= internal_cpu_0_data_master_requests_nios2_clock_4_in;
  --allow new arb cycle for nios2_clock_4/in, which is an e_assign
  nios2_clock_4_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_4_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_4_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_4_in_reset_n assignment, which is an e_assign
  nios2_clock_4_in_reset_n <= reset_n;
  --nios2_clock_4_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_4_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_4_in_begins_xfer) = '1'), nios2_clock_4_in_unreg_firsttransfer, nios2_clock_4_in_reg_firsttransfer);
  --nios2_clock_4_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_4_in_unreg_firsttransfer <= NOT ((nios2_clock_4_in_slavearbiterlockenable AND nios2_clock_4_in_any_continuerequest));
  --nios2_clock_4_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_4_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_4_in_begins_xfer) = '1' then 
        nios2_clock_4_in_reg_firsttransfer <= nios2_clock_4_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_4_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_4_in_beginbursttransfer_internal <= nios2_clock_4_in_begins_xfer;
  --nios2_clock_4_in_read assignment, which is an e_mux
  nios2_clock_4_in_read <= internal_cpu_0_data_master_granted_nios2_clock_4_in AND cpu_0_data_master_read;
  --nios2_clock_4_in_write assignment, which is an e_mux
  nios2_clock_4_in_write <= internal_cpu_0_data_master_granted_nios2_clock_4_in AND cpu_0_data_master_write;
  shifted_address_to_nios2_clock_4_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_4_in_address mux, which is an e_mux
  nios2_clock_4_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_4_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --slaveid nios2_clock_4_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_4_in_nativeaddress <= Vector_To_Std_Logic(A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")));
  --d1_nios2_clock_4_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_4_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_4_in_end_xfer <= nios2_clock_4_in_end_xfer;
    end if;

  end process;

  --nios2_clock_4_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_4_in_waits_for_read <= nios2_clock_4_in_in_a_read_cycle AND internal_nios2_clock_4_in_waitrequest_from_sa;
  --nios2_clock_4_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_4_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_4_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_4_in_in_a_read_cycle;
  --nios2_clock_4_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_4_in_waits_for_write <= nios2_clock_4_in_in_a_write_cycle AND internal_nios2_clock_4_in_waitrequest_from_sa;
  --nios2_clock_4_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_4_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_4_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_4_in_in_a_write_cycle;
  wait_for_nios2_clock_4_in_counter <= std_logic'('0');
  --nios2_clock_4_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_4_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_4_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_4_in <= internal_cpu_0_data_master_granted_nios2_clock_4_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_4_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_4_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_4_in <= internal_cpu_0_data_master_requests_nios2_clock_4_in;
  --vhdl renameroo for output signals
  nios2_clock_4_in_waitrequest_from_sa <= internal_nios2_clock_4_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_4/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_4_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_4_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_4_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_4_out_granted_sysid_control_slave : IN STD_LOGIC;
                 signal nios2_clock_4_out_qualified_request_sysid_control_slave : IN STD_LOGIC;
                 signal nios2_clock_4_out_read : IN STD_LOGIC;
                 signal nios2_clock_4_out_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                 signal nios2_clock_4_out_requests_sysid_control_slave : IN STD_LOGIC;
                 signal nios2_clock_4_out_write : IN STD_LOGIC;
                 signal nios2_clock_4_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal nios2_clock_4_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_4_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_4_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_4_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_4_out_arbitrator;


architecture europa of nios2_clock_4_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_4_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_nios2_clock_4_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_4_out_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_4_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_4_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_4_out_run :  STD_LOGIC;
                signal nios2_clock_4_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_4_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_4_out_qualified_request_sysid_control_slave OR NOT nios2_clock_4_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sysid_control_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_4_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_4_out_qualified_request_sysid_control_slave OR NOT nios2_clock_4_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_4_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_4_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_4_out_address_to_slave <= nios2_clock_4_out_address;
  --nios2_clock_4/out readdata mux, which is an e_mux
  nios2_clock_4_out_readdata <= sysid_control_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_4_out_waitrequest <= NOT nios2_clock_4_out_run;
  --nios2_clock_4_out_reset_n assignment, which is an e_assign
  nios2_clock_4_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_4_out_address_to_slave <= internal_nios2_clock_4_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_4_out_waitrequest <= internal_nios2_clock_4_out_waitrequest;
--synthesis translate_off
    --nios2_clock_4_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_4_out_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        nios2_clock_4_out_address_last_time <= nios2_clock_4_out_address;
      end if;

    end process;

    --nios2_clock_4/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_4_out_waitrequest AND ((nios2_clock_4_out_read OR nios2_clock_4_out_write));
      end if;

    end process;

    --nios2_clock_4_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line67 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_4_out_address /= nios2_clock_4_out_address_last_time))))) = '1' then 
          write(write_line67, now);
          write(write_line67, string'(": "));
          write(write_line67, string'("nios2_clock_4_out_address did not heed wait!!!"));
          write(output, write_line67.all);
          deallocate (write_line67);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_4_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_4_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_4_out_byteenable_last_time <= nios2_clock_4_out_byteenable;
      end if;

    end process;

    --nios2_clock_4_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line68 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_4_out_byteenable /= nios2_clock_4_out_byteenable_last_time))))) = '1' then 
          write(write_line68, now);
          write(write_line68, string'(": "));
          write(write_line68, string'("nios2_clock_4_out_byteenable did not heed wait!!!"));
          write(output, write_line68.all);
          deallocate (write_line68);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_4_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_4_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_4_out_read_last_time <= nios2_clock_4_out_read;
      end if;

    end process;

    --nios2_clock_4_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line69 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_4_out_read) /= std_logic'(nios2_clock_4_out_read_last_time)))))) = '1' then 
          write(write_line69, now);
          write(write_line69, string'(": "));
          write(write_line69, string'("nios2_clock_4_out_read did not heed wait!!!"));
          write(output, write_line69.all);
          deallocate (write_line69);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_4_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_4_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_4_out_write_last_time <= nios2_clock_4_out_write;
      end if;

    end process;

    --nios2_clock_4_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line70 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_4_out_write) /= std_logic'(nios2_clock_4_out_write_last_time)))))) = '1' then 
          write(write_line70, now);
          write(write_line70, string'(": "));
          write(write_line70, string'("nios2_clock_4_out_write did not heed wait!!!"));
          write(output, write_line70.all);
          deallocate (write_line70);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_4_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_4_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_4_out_writedata_last_time <= nios2_clock_4_out_writedata;
      end if;

    end process;

    --nios2_clock_4_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line71 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_4_out_writedata /= nios2_clock_4_out_writedata_last_time)))) AND nios2_clock_4_out_write)) = '1' then 
          write(write_line71, now);
          write(write_line71, string'(": "));
          write(write_line71, string'("nios2_clock_4_out_writedata did not heed wait!!!"));
          write(output, write_line71.all);
          deallocate (write_line71);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_5_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_5_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_5_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_5_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_5_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_5_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_5_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_5_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_5_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_5_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_5_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_5_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_5_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_5_in_read : OUT STD_LOGIC;
                 signal nios2_clock_5_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_5_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_5_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_5_in_write : OUT STD_LOGIC;
                 signal nios2_clock_5_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_clock_5_in_arbitrator;


architecture europa of nios2_clock_5_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_5_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_5_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_5_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_5_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_5_in :  STD_LOGIC;
                signal internal_nios2_clock_5_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_5_in_allgrants :  STD_LOGIC;
                signal nios2_clock_5_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_5_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_5_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_5_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_5_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_5_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_5_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_5_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_5_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_5_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_5_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_5_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_5_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_5_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_5_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_5_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_5_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_5_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_5_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_5_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_5_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_5_in_waits_for_write :  STD_LOGIC;
                signal wait_for_nios2_clock_5_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_5_in_end_xfer;
    end if;

  end process;

  nios2_clock_5_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_5_in);
  --assign nios2_clock_5_in_readdata_from_sa = nios2_clock_5_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_5_in_readdata_from_sa <= nios2_clock_5_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_5_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000000100000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_5_in_waitrequest_from_sa = nios2_clock_5_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_5_in_waitrequest_from_sa <= nios2_clock_5_in_waitrequest;
  --nios2_clock_5_in_arb_share_counter set values, which is an e_mux
  nios2_clock_5_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_5_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_5_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_5_in;
  --nios2_clock_5_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_5_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_5_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_5_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_5_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_5_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_5_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_5_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_5_in_allgrants all slave grants, which is an e_mux
  nios2_clock_5_in_allgrants <= nios2_clock_5_in_grant_vector;
  --nios2_clock_5_in_end_xfer assignment, which is an e_assign
  nios2_clock_5_in_end_xfer <= NOT ((nios2_clock_5_in_waits_for_read OR nios2_clock_5_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_5_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_5_in <= nios2_clock_5_in_end_xfer AND (((NOT nios2_clock_5_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_5_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_5_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_5_in AND nios2_clock_5_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_5_in AND NOT nios2_clock_5_in_non_bursting_master_requests));
  --nios2_clock_5_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_5_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_5_in_arb_counter_enable) = '1' then 
        nios2_clock_5_in_arb_share_counter <= nios2_clock_5_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_5_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_5_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_5_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_5_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_5_in AND NOT nios2_clock_5_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_5_in_slavearbiterlockenable <= or_reduce(nios2_clock_5_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_5/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_5_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_5_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_5_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_5_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_5/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_5_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_5_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_5_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_5_in <= internal_cpu_0_data_master_requests_nios2_clock_5_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_5_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_5_in <= (internal_cpu_0_data_master_granted_nios2_clock_5_in AND cpu_0_data_master_read) AND NOT nios2_clock_5_in_waits_for_read;
  --nios2_clock_5_in_writedata mux, which is an e_mux
  nios2_clock_5_in_writedata <= cpu_0_data_master_writedata;
  --assign nios2_clock_5_in_endofpacket_from_sa = nios2_clock_5_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_5_in_endofpacket_from_sa <= nios2_clock_5_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_5_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_5_in;
  --cpu_0/data_master saved-grant nios2_clock_5/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_5_in <= internal_cpu_0_data_master_requests_nios2_clock_5_in;
  --allow new arb cycle for nios2_clock_5/in, which is an e_assign
  nios2_clock_5_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_5_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_5_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_5_in_reset_n assignment, which is an e_assign
  nios2_clock_5_in_reset_n <= reset_n;
  --nios2_clock_5_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_5_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_5_in_begins_xfer) = '1'), nios2_clock_5_in_unreg_firsttransfer, nios2_clock_5_in_reg_firsttransfer);
  --nios2_clock_5_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_5_in_unreg_firsttransfer <= NOT ((nios2_clock_5_in_slavearbiterlockenable AND nios2_clock_5_in_any_continuerequest));
  --nios2_clock_5_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_5_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_5_in_begins_xfer) = '1' then 
        nios2_clock_5_in_reg_firsttransfer <= nios2_clock_5_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_5_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_5_in_beginbursttransfer_internal <= nios2_clock_5_in_begins_xfer;
  --nios2_clock_5_in_read assignment, which is an e_mux
  nios2_clock_5_in_read <= internal_cpu_0_data_master_granted_nios2_clock_5_in AND cpu_0_data_master_read;
  --nios2_clock_5_in_write assignment, which is an e_mux
  nios2_clock_5_in_write <= internal_cpu_0_data_master_granted_nios2_clock_5_in AND cpu_0_data_master_write;
  --nios2_clock_5_in_address mux, which is an e_mux
  nios2_clock_5_in_address <= cpu_0_data_master_address_to_slave (3 DOWNTO 0);
  --slaveid nios2_clock_5_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_5_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_5_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_5_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_5_in_end_xfer <= nios2_clock_5_in_end_xfer;
    end if;

  end process;

  --nios2_clock_5_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_5_in_waits_for_read <= nios2_clock_5_in_in_a_read_cycle AND internal_nios2_clock_5_in_waitrequest_from_sa;
  --nios2_clock_5_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_5_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_5_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_5_in_in_a_read_cycle;
  --nios2_clock_5_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_5_in_waits_for_write <= nios2_clock_5_in_in_a_write_cycle AND internal_nios2_clock_5_in_waitrequest_from_sa;
  --nios2_clock_5_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_5_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_5_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_5_in_in_a_write_cycle;
  wait_for_nios2_clock_5_in_counter <= std_logic'('0');
  --nios2_clock_5_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_5_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_5_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_5_in <= internal_cpu_0_data_master_granted_nios2_clock_5_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_5_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_5_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_5_in <= internal_cpu_0_data_master_requests_nios2_clock_5_in;
  --vhdl renameroo for output signals
  nios2_clock_5_in_waitrequest_from_sa <= internal_nios2_clock_5_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_5/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_5_out_arbitrator is 
        port (
              -- inputs:
                 signal altpll_0_pll_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_altpll_0_pll_slave_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_5_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_5_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_5_out_granted_altpll_0_pll_slave : IN STD_LOGIC;
                 signal nios2_clock_5_out_qualified_request_altpll_0_pll_slave : IN STD_LOGIC;
                 signal nios2_clock_5_out_read : IN STD_LOGIC;
                 signal nios2_clock_5_out_read_data_valid_altpll_0_pll_slave : IN STD_LOGIC;
                 signal nios2_clock_5_out_requests_altpll_0_pll_slave : IN STD_LOGIC;
                 signal nios2_clock_5_out_write : IN STD_LOGIC;
                 signal nios2_clock_5_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_5_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_5_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_5_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_5_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_5_out_arbitrator;


architecture europa of nios2_clock_5_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_5_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_clock_5_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_5_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_5_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_5_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_5_out_run :  STD_LOGIC;
                signal nios2_clock_5_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_5_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_5_out_qualified_request_altpll_0_pll_slave OR NOT ((nios2_clock_5_out_read OR nios2_clock_5_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_5_out_read OR nios2_clock_5_out_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_5_out_qualified_request_altpll_0_pll_slave OR NOT ((nios2_clock_5_out_read OR nios2_clock_5_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_5_out_read OR nios2_clock_5_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_5_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_5_out_address_to_slave <= nios2_clock_5_out_address;
  --nios2_clock_5/out readdata mux, which is an e_mux
  nios2_clock_5_out_readdata <= altpll_0_pll_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_5_out_waitrequest <= NOT nios2_clock_5_out_run;
  --nios2_clock_5_out_reset_n assignment, which is an e_assign
  nios2_clock_5_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_5_out_address_to_slave <= internal_nios2_clock_5_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_5_out_waitrequest <= internal_nios2_clock_5_out_waitrequest;
--synthesis translate_off
    --nios2_clock_5_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_5_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_5_out_address_last_time <= nios2_clock_5_out_address;
      end if;

    end process;

    --nios2_clock_5/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_5_out_waitrequest AND ((nios2_clock_5_out_read OR nios2_clock_5_out_write));
      end if;

    end process;

    --nios2_clock_5_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line72 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_5_out_address /= nios2_clock_5_out_address_last_time))))) = '1' then 
          write(write_line72, now);
          write(write_line72, string'(": "));
          write(write_line72, string'("nios2_clock_5_out_address did not heed wait!!!"));
          write(output, write_line72.all);
          deallocate (write_line72);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_5_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_5_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_5_out_byteenable_last_time <= nios2_clock_5_out_byteenable;
      end if;

    end process;

    --nios2_clock_5_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line73 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_5_out_byteenable /= nios2_clock_5_out_byteenable_last_time))))) = '1' then 
          write(write_line73, now);
          write(write_line73, string'(": "));
          write(write_line73, string'("nios2_clock_5_out_byteenable did not heed wait!!!"));
          write(output, write_line73.all);
          deallocate (write_line73);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_5_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_5_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_5_out_read_last_time <= nios2_clock_5_out_read;
      end if;

    end process;

    --nios2_clock_5_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line74 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_5_out_read) /= std_logic'(nios2_clock_5_out_read_last_time)))))) = '1' then 
          write(write_line74, now);
          write(write_line74, string'(": "));
          write(write_line74, string'("nios2_clock_5_out_read did not heed wait!!!"));
          write(output, write_line74.all);
          deallocate (write_line74);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_5_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_5_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_5_out_write_last_time <= nios2_clock_5_out_write;
      end if;

    end process;

    --nios2_clock_5_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line75 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_5_out_write) /= std_logic'(nios2_clock_5_out_write_last_time)))))) = '1' then 
          write(write_line75, now);
          write(write_line75, string'(": "));
          write(write_line75, string'("nios2_clock_5_out_write did not heed wait!!!"));
          write(output, write_line75.all);
          deallocate (write_line75);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_5_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_5_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_5_out_writedata_last_time <= nios2_clock_5_out_writedata;
      end if;

    end process;

    --nios2_clock_5_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line76 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_5_out_writedata /= nios2_clock_5_out_writedata_last_time)))) AND nios2_clock_5_out_write)) = '1' then 
          write(write_line76, now);
          write(write_line76, string'(": "));
          write(write_line76, string'("nios2_clock_5_out_writedata did not heed wait!!!"));
          write(output, write_line76.all);
          deallocate (write_line76);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_6_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_6_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_6_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_6_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_6_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_6_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_6_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_6_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_6_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_6_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_6_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_6_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_6_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_6_in_read : OUT STD_LOGIC;
                 signal nios2_clock_6_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_6_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_6_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_6_in_write : OUT STD_LOGIC;
                 signal nios2_clock_6_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_clock_6_in_arbitrator;


architecture europa of nios2_clock_6_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_6_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_6_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_6_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_6_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_6_in :  STD_LOGIC;
                signal internal_nios2_clock_6_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_6_in_allgrants :  STD_LOGIC;
                signal nios2_clock_6_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_6_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_6_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_6_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_6_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_6_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_6_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_6_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_6_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_6_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_6_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_6_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_6_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_6_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_6_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_6_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_6_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_6_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_6_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_6_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_6_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_6_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_6_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_6_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_6_in_end_xfer;
    end if;

  end process;

  nios2_clock_6_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_6_in);
  --assign nios2_clock_6_in_readdata_from_sa = nios2_clock_6_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_6_in_readdata_from_sa <= nios2_clock_6_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_6_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000000110000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_6_in_waitrequest_from_sa = nios2_clock_6_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_6_in_waitrequest_from_sa <= nios2_clock_6_in_waitrequest;
  --nios2_clock_6_in_arb_share_counter set values, which is an e_mux
  nios2_clock_6_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_6_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_6_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_6_in;
  --nios2_clock_6_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_6_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_6_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_6_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_6_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_6_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_6_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_6_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_6_in_allgrants all slave grants, which is an e_mux
  nios2_clock_6_in_allgrants <= nios2_clock_6_in_grant_vector;
  --nios2_clock_6_in_end_xfer assignment, which is an e_assign
  nios2_clock_6_in_end_xfer <= NOT ((nios2_clock_6_in_waits_for_read OR nios2_clock_6_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_6_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_6_in <= nios2_clock_6_in_end_xfer AND (((NOT nios2_clock_6_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_6_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_6_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_6_in AND nios2_clock_6_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_6_in AND NOT nios2_clock_6_in_non_bursting_master_requests));
  --nios2_clock_6_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_6_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_6_in_arb_counter_enable) = '1' then 
        nios2_clock_6_in_arb_share_counter <= nios2_clock_6_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_6_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_6_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_6_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_6_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_6_in AND NOT nios2_clock_6_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_6_in_slavearbiterlockenable <= or_reduce(nios2_clock_6_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_6/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_6_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_6_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_6_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_6_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_6/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_6_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_6_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_6_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_6_in <= internal_cpu_0_data_master_requests_nios2_clock_6_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_6_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_6_in <= (internal_cpu_0_data_master_granted_nios2_clock_6_in AND cpu_0_data_master_read) AND NOT nios2_clock_6_in_waits_for_read;
  --nios2_clock_6_in_writedata mux, which is an e_mux
  nios2_clock_6_in_writedata <= cpu_0_data_master_writedata;
  --assign nios2_clock_6_in_endofpacket_from_sa = nios2_clock_6_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_6_in_endofpacket_from_sa <= nios2_clock_6_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_6_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_6_in;
  --cpu_0/data_master saved-grant nios2_clock_6/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_6_in <= internal_cpu_0_data_master_requests_nios2_clock_6_in;
  --allow new arb cycle for nios2_clock_6/in, which is an e_assign
  nios2_clock_6_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_6_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_6_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_6_in_reset_n assignment, which is an e_assign
  nios2_clock_6_in_reset_n <= reset_n;
  --nios2_clock_6_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_6_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_6_in_begins_xfer) = '1'), nios2_clock_6_in_unreg_firsttransfer, nios2_clock_6_in_reg_firsttransfer);
  --nios2_clock_6_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_6_in_unreg_firsttransfer <= NOT ((nios2_clock_6_in_slavearbiterlockenable AND nios2_clock_6_in_any_continuerequest));
  --nios2_clock_6_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_6_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_6_in_begins_xfer) = '1' then 
        nios2_clock_6_in_reg_firsttransfer <= nios2_clock_6_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_6_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_6_in_beginbursttransfer_internal <= nios2_clock_6_in_begins_xfer;
  --nios2_clock_6_in_read assignment, which is an e_mux
  nios2_clock_6_in_read <= internal_cpu_0_data_master_granted_nios2_clock_6_in AND cpu_0_data_master_read;
  --nios2_clock_6_in_write assignment, which is an e_mux
  nios2_clock_6_in_write <= internal_cpu_0_data_master_granted_nios2_clock_6_in AND cpu_0_data_master_write;
  shifted_address_to_nios2_clock_6_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_6_in_address mux, which is an e_mux
  nios2_clock_6_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_6_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --slaveid nios2_clock_6_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_6_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_6_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_6_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_6_in_end_xfer <= nios2_clock_6_in_end_xfer;
    end if;

  end process;

  --nios2_clock_6_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_6_in_waits_for_read <= nios2_clock_6_in_in_a_read_cycle AND internal_nios2_clock_6_in_waitrequest_from_sa;
  --nios2_clock_6_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_6_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_6_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_6_in_in_a_read_cycle;
  --nios2_clock_6_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_6_in_waits_for_write <= nios2_clock_6_in_in_a_write_cycle AND internal_nios2_clock_6_in_waitrequest_from_sa;
  --nios2_clock_6_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_6_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_6_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_6_in_in_a_write_cycle;
  wait_for_nios2_clock_6_in_counter <= std_logic'('0');
  --nios2_clock_6_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_6_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_6_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_6_in <= internal_cpu_0_data_master_granted_nios2_clock_6_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_6_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_6_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_6_in <= internal_cpu_0_data_master_requests_nios2_clock_6_in;
  --vhdl renameroo for output signals
  nios2_clock_6_in_waitrequest_from_sa <= internal_nios2_clock_6_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_6/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_6_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_gen_code_value_pio_0_s1_end_xfer : IN STD_LOGIC;
                 signal gen_code_value_pio_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal nios2_clock_6_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_6_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_6_out_granted_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_6_out_read : IN STD_LOGIC;
                 signal nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_6_out_requests_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_6_out_write : IN STD_LOGIC;
                 signal nios2_clock_6_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_6_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_6_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_6_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_6_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_6_out_arbitrator;


architecture europa of nios2_clock_6_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_6_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_clock_6_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_6_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_6_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_6_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_6_out_run :  STD_LOGIC;
                signal nios2_clock_6_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_6_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 OR NOT nios2_clock_6_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_gen_code_value_pio_0_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_6_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 OR NOT nios2_clock_6_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_6_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_6_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_6_out_address_to_slave <= nios2_clock_6_out_address;
  --nios2_clock_6/out readdata mux, which is an e_mux
  nios2_clock_6_out_readdata <= std_logic_vector'("00000000") & (gen_code_value_pio_0_s1_readdata_from_sa);
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_6_out_waitrequest <= NOT nios2_clock_6_out_run;
  --nios2_clock_6_out_reset_n assignment, which is an e_assign
  nios2_clock_6_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_6_out_address_to_slave <= internal_nios2_clock_6_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_6_out_waitrequest <= internal_nios2_clock_6_out_waitrequest;
--synthesis translate_off
    --nios2_clock_6_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_6_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_6_out_address_last_time <= nios2_clock_6_out_address;
      end if;

    end process;

    --nios2_clock_6/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_6_out_waitrequest AND ((nios2_clock_6_out_read OR nios2_clock_6_out_write));
      end if;

    end process;

    --nios2_clock_6_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line77 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_6_out_address /= nios2_clock_6_out_address_last_time))))) = '1' then 
          write(write_line77, now);
          write(write_line77, string'(": "));
          write(write_line77, string'("nios2_clock_6_out_address did not heed wait!!!"));
          write(output, write_line77.all);
          deallocate (write_line77);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_6_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_6_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_6_out_byteenable_last_time <= nios2_clock_6_out_byteenable;
      end if;

    end process;

    --nios2_clock_6_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line78 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_6_out_byteenable /= nios2_clock_6_out_byteenable_last_time))))) = '1' then 
          write(write_line78, now);
          write(write_line78, string'(": "));
          write(write_line78, string'("nios2_clock_6_out_byteenable did not heed wait!!!"));
          write(output, write_line78.all);
          deallocate (write_line78);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_6_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_6_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_6_out_read_last_time <= nios2_clock_6_out_read;
      end if;

    end process;

    --nios2_clock_6_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line79 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_6_out_read) /= std_logic'(nios2_clock_6_out_read_last_time)))))) = '1' then 
          write(write_line79, now);
          write(write_line79, string'(": "));
          write(write_line79, string'("nios2_clock_6_out_read did not heed wait!!!"));
          write(output, write_line79.all);
          deallocate (write_line79);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_6_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_6_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_6_out_write_last_time <= nios2_clock_6_out_write;
      end if;

    end process;

    --nios2_clock_6_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line80 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_6_out_write) /= std_logic'(nios2_clock_6_out_write_last_time)))))) = '1' then 
          write(write_line80, now);
          write(write_line80, string'(": "));
          write(write_line80, string'("nios2_clock_6_out_write did not heed wait!!!"));
          write(output, write_line80.all);
          deallocate (write_line80);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_6_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_6_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_6_out_writedata_last_time <= nios2_clock_6_out_writedata;
      end if;

    end process;

    --nios2_clock_6_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line81 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_6_out_writedata /= nios2_clock_6_out_writedata_last_time)))) AND nios2_clock_6_out_write)) = '1' then 
          write(write_line81, now);
          write(write_line81, string'(": "));
          write(write_line81, string'("nios2_clock_6_out_writedata did not heed wait!!!"));
          write(output, write_line81.all);
          deallocate (write_line81);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_7_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_7_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_7_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_7_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_nios2_clock_7_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_7_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_7_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_7_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_7_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_7_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_7_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_7_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_7_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_7_in_read : OUT STD_LOGIC;
                 signal nios2_clock_7_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_7_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_7_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_7_in_write : OUT STD_LOGIC;
                 signal nios2_clock_7_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_clock_7_in_arbitrator;


architecture europa of nios2_clock_7_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_7_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_7_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_nios2_clock_7_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_7_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_7_in :  STD_LOGIC;
                signal internal_nios2_clock_7_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_7_in_allgrants :  STD_LOGIC;
                signal nios2_clock_7_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_7_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_7_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_7_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_7_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_7_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_7_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_7_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_7_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_7_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_7_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_7_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_7_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_7_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_7_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_7_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_7_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_7_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_7_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_7_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_7_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_7_in_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_nios2_clock_7_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_nios2_clock_7_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_7_in_end_xfer;
    end if;

  end process;

  nios2_clock_7_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_7_in);
  --assign nios2_clock_7_in_readdata_from_sa = nios2_clock_7_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_7_in_readdata_from_sa <= nios2_clock_7_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_7_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000010001000001000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_7_in_waitrequest_from_sa = nios2_clock_7_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_7_in_waitrequest_from_sa <= nios2_clock_7_in_waitrequest;
  --nios2_clock_7_in_arb_share_counter set values, which is an e_mux
  nios2_clock_7_in_arb_share_set_values <= std_logic_vector'("01");
  --nios2_clock_7_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_7_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_7_in;
  --nios2_clock_7_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_7_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_7_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_7_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_7_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_7_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_7_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_7_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_7_in_allgrants all slave grants, which is an e_mux
  nios2_clock_7_in_allgrants <= nios2_clock_7_in_grant_vector;
  --nios2_clock_7_in_end_xfer assignment, which is an e_assign
  nios2_clock_7_in_end_xfer <= NOT ((nios2_clock_7_in_waits_for_read OR nios2_clock_7_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_7_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_7_in <= nios2_clock_7_in_end_xfer AND (((NOT nios2_clock_7_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_7_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_7_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_7_in AND nios2_clock_7_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_7_in AND NOT nios2_clock_7_in_non_bursting_master_requests));
  --nios2_clock_7_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_7_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_7_in_arb_counter_enable) = '1' then 
        nios2_clock_7_in_arb_share_counter <= nios2_clock_7_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_7_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_7_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_7_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_7_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_7_in AND NOT nios2_clock_7_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_7_in_slavearbiterlockenable <= or_reduce(nios2_clock_7_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_7/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_7_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_7_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_7_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_7_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_7/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_7_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_7_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_7_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_7_in <= internal_cpu_0_data_master_requests_nios2_clock_7_in AND NOT ((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_7_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_7_in <= (internal_cpu_0_data_master_granted_nios2_clock_7_in AND cpu_0_data_master_read) AND NOT nios2_clock_7_in_waits_for_read;
  --nios2_clock_7_in_writedata mux, which is an e_mux
  nios2_clock_7_in_writedata <= cpu_0_data_master_writedata;
  --assign nios2_clock_7_in_endofpacket_from_sa = nios2_clock_7_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_7_in_endofpacket_from_sa <= nios2_clock_7_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_7_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_7_in;
  --cpu_0/data_master saved-grant nios2_clock_7/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_7_in <= internal_cpu_0_data_master_requests_nios2_clock_7_in;
  --allow new arb cycle for nios2_clock_7/in, which is an e_assign
  nios2_clock_7_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_7_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_7_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_7_in_reset_n assignment, which is an e_assign
  nios2_clock_7_in_reset_n <= reset_n;
  --nios2_clock_7_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_7_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_7_in_begins_xfer) = '1'), nios2_clock_7_in_unreg_firsttransfer, nios2_clock_7_in_reg_firsttransfer);
  --nios2_clock_7_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_7_in_unreg_firsttransfer <= NOT ((nios2_clock_7_in_slavearbiterlockenable AND nios2_clock_7_in_any_continuerequest));
  --nios2_clock_7_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_7_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_7_in_begins_xfer) = '1' then 
        nios2_clock_7_in_reg_firsttransfer <= nios2_clock_7_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_7_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_7_in_beginbursttransfer_internal <= nios2_clock_7_in_begins_xfer;
  --nios2_clock_7_in_read assignment, which is an e_mux
  nios2_clock_7_in_read <= internal_cpu_0_data_master_granted_nios2_clock_7_in AND cpu_0_data_master_read;
  --nios2_clock_7_in_write assignment, which is an e_mux
  nios2_clock_7_in_write <= internal_cpu_0_data_master_granted_nios2_clock_7_in AND cpu_0_data_master_write;
  shifted_address_to_nios2_clock_7_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --nios2_clock_7_in_address mux, which is an e_mux
  nios2_clock_7_in_address <= A_EXT (A_SRL(shifted_address_to_nios2_clock_7_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --slaveid nios2_clock_7_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_7_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_nios2_clock_7_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_7_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_7_in_end_xfer <= nios2_clock_7_in_end_xfer;
    end if;

  end process;

  --nios2_clock_7_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_7_in_waits_for_read <= nios2_clock_7_in_in_a_read_cycle AND internal_nios2_clock_7_in_waitrequest_from_sa;
  --nios2_clock_7_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_7_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_7_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_7_in_in_a_read_cycle;
  --nios2_clock_7_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_7_in_waits_for_write <= nios2_clock_7_in_in_a_write_cycle AND internal_nios2_clock_7_in_waitrequest_from_sa;
  --nios2_clock_7_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_7_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_7_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_7_in_in_a_write_cycle;
  wait_for_nios2_clock_7_in_counter <= std_logic'('0');
  --nios2_clock_7_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_7_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_7_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_7_in <= internal_cpu_0_data_master_granted_nios2_clock_7_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_7_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_7_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_7_in <= internal_cpu_0_data_master_requests_nios2_clock_7_in;
  --vhdl renameroo for output signals
  nios2_clock_7_in_waitrequest_from_sa <= internal_nios2_clock_7_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_7/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_7_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_gen_code_value_pio_1_s1_end_xfer : IN STD_LOGIC;
                 signal gen_code_value_pio_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal nios2_clock_7_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_7_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_7_out_granted_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                 signal nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                 signal nios2_clock_7_out_read : IN STD_LOGIC;
                 signal nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                 signal nios2_clock_7_out_requests_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                 signal nios2_clock_7_out_write : IN STD_LOGIC;
                 signal nios2_clock_7_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_7_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_7_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_7_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_7_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_7_out_arbitrator;


architecture europa of nios2_clock_7_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_7_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_clock_7_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_7_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_7_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_7_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_7_out_run :  STD_LOGIC;
                signal nios2_clock_7_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_7_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 OR NOT nios2_clock_7_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_gen_code_value_pio_1_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_7_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 OR NOT nios2_clock_7_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_7_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_7_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_7_out_address_to_slave <= nios2_clock_7_out_address;
  --nios2_clock_7/out readdata mux, which is an e_mux
  nios2_clock_7_out_readdata <= std_logic_vector'("00000000") & (gen_code_value_pio_1_s1_readdata_from_sa);
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_7_out_waitrequest <= NOT nios2_clock_7_out_run;
  --nios2_clock_7_out_reset_n assignment, which is an e_assign
  nios2_clock_7_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_7_out_address_to_slave <= internal_nios2_clock_7_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_7_out_waitrequest <= internal_nios2_clock_7_out_waitrequest;
--synthesis translate_off
    --nios2_clock_7_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_7_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_7_out_address_last_time <= nios2_clock_7_out_address;
      end if;

    end process;

    --nios2_clock_7/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_7_out_waitrequest AND ((nios2_clock_7_out_read OR nios2_clock_7_out_write));
      end if;

    end process;

    --nios2_clock_7_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line82 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_7_out_address /= nios2_clock_7_out_address_last_time))))) = '1' then 
          write(write_line82, now);
          write(write_line82, string'(": "));
          write(write_line82, string'("nios2_clock_7_out_address did not heed wait!!!"));
          write(output, write_line82.all);
          deallocate (write_line82);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_7_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_7_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_clock_7_out_byteenable_last_time <= nios2_clock_7_out_byteenable;
      end if;

    end process;

    --nios2_clock_7_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line83 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_7_out_byteenable /= nios2_clock_7_out_byteenable_last_time))))) = '1' then 
          write(write_line83, now);
          write(write_line83, string'(": "));
          write(write_line83, string'("nios2_clock_7_out_byteenable did not heed wait!!!"));
          write(output, write_line83.all);
          deallocate (write_line83);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_7_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_7_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_7_out_read_last_time <= nios2_clock_7_out_read;
      end if;

    end process;

    --nios2_clock_7_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line84 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_7_out_read) /= std_logic'(nios2_clock_7_out_read_last_time)))))) = '1' then 
          write(write_line84, now);
          write(write_line84, string'(": "));
          write(write_line84, string'("nios2_clock_7_out_read did not heed wait!!!"));
          write(output, write_line84.all);
          deallocate (write_line84);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_7_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_7_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_7_out_write_last_time <= nios2_clock_7_out_write;
      end if;

    end process;

    --nios2_clock_7_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line85 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_7_out_write) /= std_logic'(nios2_clock_7_out_write_last_time)))))) = '1' then 
          write(write_line85, now);
          write(write_line85, string'(": "));
          write(write_line85, string'("nios2_clock_7_out_write did not heed wait!!!"));
          write(output, write_line85.all);
          deallocate (write_line85);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_7_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_7_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_7_out_writedata_last_time <= nios2_clock_7_out_writedata;
      end if;

    end process;

    --nios2_clock_7_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line86 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_7_out_writedata /= nios2_clock_7_out_writedata_last_time)))) AND nios2_clock_7_out_write)) = '1' then 
          write(write_line86, now);
          write(write_line86, string'(": "));
          write(write_line86, string'("nios2_clock_7_out_writedata did not heed wait!!!"));
          write(output, write_line86.all);
          deallocate (write_line86);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_8_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_0_instruction_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal nios2_clock_8_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_8_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_8_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_instruction_master_granted_nios2_clock_8_in : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_nios2_clock_8_in : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_nios2_clock_8_in : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_nios2_clock_8_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_8_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_8_in_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_8_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_8_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_8_in_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal nios2_clock_8_in_read : OUT STD_LOGIC;
                 signal nios2_clock_8_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_8_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_8_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_8_in_write : OUT STD_LOGIC
              );
end entity nios2_clock_8_in_arbitrator;


architecture europa of nios2_clock_8_in_arbitrator is
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_nios2_clock_8_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_8_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_nios2_clock_8_in :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_nios2_clock_8_in :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_nios2_clock_8_in :  STD_LOGIC;
                signal internal_nios2_clock_8_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_8_in_allgrants :  STD_LOGIC;
                signal nios2_clock_8_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_8_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_8_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_8_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_8_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_8_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_8_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_8_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_8_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_8_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_8_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_8_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_8_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_8_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_8_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_8_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_8_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_8_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_8_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_8_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_8_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_8_in_waits_for_write :  STD_LOGIC;
                signal wait_for_nios2_clock_8_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_8_in_end_xfer;
    end if;

  end process;

  nios2_clock_8_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_instruction_master_qualified_request_nios2_clock_8_in);
  --assign nios2_clock_8_in_readdata_from_sa = nios2_clock_8_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_8_in_readdata_from_sa <= nios2_clock_8_in_readdata;
  internal_cpu_0_instruction_master_requests_nios2_clock_8_in <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(24 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("0100000000000000000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --assign nios2_clock_8_in_waitrequest_from_sa = nios2_clock_8_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_8_in_waitrequest_from_sa <= nios2_clock_8_in_waitrequest;
  --nios2_clock_8_in_arb_share_counter set values, which is an e_mux
  nios2_clock_8_in_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_instruction_master_granted_nios2_clock_8_in)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001")), 2);
  --nios2_clock_8_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_8_in_non_bursting_master_requests <= internal_cpu_0_instruction_master_requests_nios2_clock_8_in;
  --nios2_clock_8_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_8_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_8_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_8_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_8_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_8_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_8_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_8_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_8_in_allgrants all slave grants, which is an e_mux
  nios2_clock_8_in_allgrants <= nios2_clock_8_in_grant_vector;
  --nios2_clock_8_in_end_xfer assignment, which is an e_assign
  nios2_clock_8_in_end_xfer <= NOT ((nios2_clock_8_in_waits_for_read OR nios2_clock_8_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_8_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_8_in <= nios2_clock_8_in_end_xfer AND (((NOT nios2_clock_8_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_8_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_8_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_8_in AND nios2_clock_8_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_8_in AND NOT nios2_clock_8_in_non_bursting_master_requests));
  --nios2_clock_8_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_8_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_8_in_arb_counter_enable) = '1' then 
        nios2_clock_8_in_arb_share_counter <= nios2_clock_8_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_8_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_8_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_8_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_8_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_8_in AND NOT nios2_clock_8_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_8_in_slavearbiterlockenable <= or_reduce(nios2_clock_8_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/instruction_master nios2_clock_8/in arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= nios2_clock_8_in_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --nios2_clock_8_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_8_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_8_in_arb_share_counter_next_value);
  --cpu_0/instruction_master nios2_clock_8/in arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= nios2_clock_8_in_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --nios2_clock_8_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_8_in_any_continuerequest <= std_logic'('1');
  --cpu_0_instruction_master_continuerequest continued request, which is an e_assign
  cpu_0_instruction_master_continuerequest <= std_logic'('1');
  internal_cpu_0_instruction_master_qualified_request_nios2_clock_8_in <= internal_cpu_0_instruction_master_requests_nios2_clock_8_in AND NOT ((cpu_0_instruction_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid cpu_0_instruction_master_read_data_valid_nios2_clock_8_in, which is an e_mux
  cpu_0_instruction_master_read_data_valid_nios2_clock_8_in <= (internal_cpu_0_instruction_master_granted_nios2_clock_8_in AND cpu_0_instruction_master_read) AND NOT nios2_clock_8_in_waits_for_read;
  --assign nios2_clock_8_in_endofpacket_from_sa = nios2_clock_8_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_8_in_endofpacket_from_sa <= nios2_clock_8_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_instruction_master_granted_nios2_clock_8_in <= internal_cpu_0_instruction_master_qualified_request_nios2_clock_8_in;
  --cpu_0/instruction_master saved-grant nios2_clock_8/in, which is an e_assign
  cpu_0_instruction_master_saved_grant_nios2_clock_8_in <= internal_cpu_0_instruction_master_requests_nios2_clock_8_in;
  --allow new arb cycle for nios2_clock_8/in, which is an e_assign
  nios2_clock_8_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_8_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_8_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_8_in_reset_n assignment, which is an e_assign
  nios2_clock_8_in_reset_n <= reset_n;
  --nios2_clock_8_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_8_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_8_in_begins_xfer) = '1'), nios2_clock_8_in_unreg_firsttransfer, nios2_clock_8_in_reg_firsttransfer);
  --nios2_clock_8_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_8_in_unreg_firsttransfer <= NOT ((nios2_clock_8_in_slavearbiterlockenable AND nios2_clock_8_in_any_continuerequest));
  --nios2_clock_8_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_8_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_8_in_begins_xfer) = '1' then 
        nios2_clock_8_in_reg_firsttransfer <= nios2_clock_8_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_8_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_8_in_beginbursttransfer_internal <= nios2_clock_8_in_begins_xfer;
  --nios2_clock_8_in_read assignment, which is an e_mux
  nios2_clock_8_in_read <= internal_cpu_0_instruction_master_granted_nios2_clock_8_in AND cpu_0_instruction_master_read;
  --nios2_clock_8_in_write assignment, which is an e_mux
  nios2_clock_8_in_write <= std_logic'('0');
  --nios2_clock_8_in_address mux, which is an e_mux
  nios2_clock_8_in_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_0_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_0_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 23);
  --slaveid nios2_clock_8_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_8_in_nativeaddress <= A_EXT (A_SRL(cpu_0_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 22);
  --d1_nios2_clock_8_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_8_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_8_in_end_xfer <= nios2_clock_8_in_end_xfer;
    end if;

  end process;

  --nios2_clock_8_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_8_in_waits_for_read <= nios2_clock_8_in_in_a_read_cycle AND internal_nios2_clock_8_in_waitrequest_from_sa;
  --nios2_clock_8_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_8_in_in_a_read_cycle <= internal_cpu_0_instruction_master_granted_nios2_clock_8_in AND cpu_0_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_8_in_in_a_read_cycle;
  --nios2_clock_8_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_8_in_waits_for_write <= nios2_clock_8_in_in_a_write_cycle AND internal_nios2_clock_8_in_waitrequest_from_sa;
  --nios2_clock_8_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_8_in_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_8_in_in_a_write_cycle;
  wait_for_nios2_clock_8_in_counter <= std_logic'('0');
  --nios2_clock_8_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_8_in_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 2);
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_nios2_clock_8_in <= internal_cpu_0_instruction_master_granted_nios2_clock_8_in;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_nios2_clock_8_in <= internal_cpu_0_instruction_master_qualified_request_nios2_clock_8_in;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_nios2_clock_8_in <= internal_cpu_0_instruction_master_requests_nios2_clock_8_in;
  --vhdl renameroo for output signals
  nios2_clock_8_in_waitrequest_from_sa <= internal_nios2_clock_8_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_8/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_8_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_8_out_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_8_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_8_out_granted_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_8_out_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_8_out_read : IN STD_LOGIC;
                 signal nios2_clock_8_out_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal nios2_clock_8_out_requests_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_8_out_write : IN STD_LOGIC;
                 signal nios2_clock_8_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_8_out_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_8_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_8_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_8_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_8_out_arbitrator;


architecture europa of nios2_clock_8_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_8_out_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal internal_nios2_clock_8_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_8_out_address_last_time :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_8_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_8_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_8_out_run :  STD_LOGIC;
                signal nios2_clock_8_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_8_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((nios2_clock_8_out_qualified_request_sdram_0_s1 OR nios2_clock_8_out_read_data_valid_sdram_0_s1) OR NOT nios2_clock_8_out_requests_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_8_out_granted_sdram_0_s1 OR NOT nios2_clock_8_out_qualified_request_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT nios2_clock_8_out_qualified_request_sdram_0_s1 OR NOT nios2_clock_8_out_read) OR ((nios2_clock_8_out_read_data_valid_sdram_0_s1 AND nios2_clock_8_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_8_out_qualified_request_sdram_0_s1 OR NOT ((nios2_clock_8_out_read OR nios2_clock_8_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_0_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_8_out_read OR nios2_clock_8_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_8_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_8_out_address_to_slave <= nios2_clock_8_out_address;
  --nios2_clock_8/out readdata mux, which is an e_mux
  nios2_clock_8_out_readdata <= sdram_0_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_8_out_waitrequest <= NOT nios2_clock_8_out_run;
  --nios2_clock_8_out_reset_n assignment, which is an e_assign
  nios2_clock_8_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_8_out_address_to_slave <= internal_nios2_clock_8_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_8_out_waitrequest <= internal_nios2_clock_8_out_waitrequest;
--synthesis translate_off
    --nios2_clock_8_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_8_out_address_last_time <= std_logic_vector'("00000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_8_out_address_last_time <= nios2_clock_8_out_address;
      end if;

    end process;

    --nios2_clock_8/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_8_out_waitrequest AND ((nios2_clock_8_out_read OR nios2_clock_8_out_write));
      end if;

    end process;

    --nios2_clock_8_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line87 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_8_out_address /= nios2_clock_8_out_address_last_time))))) = '1' then 
          write(write_line87, now);
          write(write_line87, string'(": "));
          write(write_line87, string'("nios2_clock_8_out_address did not heed wait!!!"));
          write(output, write_line87.all);
          deallocate (write_line87);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_8_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_8_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_8_out_byteenable_last_time <= nios2_clock_8_out_byteenable;
      end if;

    end process;

    --nios2_clock_8_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line88 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_8_out_byteenable /= nios2_clock_8_out_byteenable_last_time))))) = '1' then 
          write(write_line88, now);
          write(write_line88, string'(": "));
          write(write_line88, string'("nios2_clock_8_out_byteenable did not heed wait!!!"));
          write(output, write_line88.all);
          deallocate (write_line88);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_8_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_8_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_8_out_read_last_time <= nios2_clock_8_out_read;
      end if;

    end process;

    --nios2_clock_8_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line89 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_8_out_read) /= std_logic'(nios2_clock_8_out_read_last_time)))))) = '1' then 
          write(write_line89, now);
          write(write_line89, string'(": "));
          write(write_line89, string'("nios2_clock_8_out_read did not heed wait!!!"));
          write(output, write_line89.all);
          deallocate (write_line89);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_8_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_8_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_8_out_write_last_time <= nios2_clock_8_out_write;
      end if;

    end process;

    --nios2_clock_8_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line90 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_8_out_write) /= std_logic'(nios2_clock_8_out_write_last_time)))))) = '1' then 
          write(write_line90, now);
          write(write_line90, string'(": "));
          write(write_line90, string'("nios2_clock_8_out_write did not heed wait!!!"));
          write(output, write_line90.all);
          deallocate (write_line90);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_8_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_8_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_8_out_writedata_last_time <= nios2_clock_8_out_writedata;
      end if;

    end process;

    --nios2_clock_8_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line91 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_8_out_writedata /= nios2_clock_8_out_writedata_last_time)))) AND nios2_clock_8_out_write)) = '1' then 
          write(write_line91, now);
          write(write_line91, string'(": "));
          write(write_line91, string'("nios2_clock_8_out_writedata did not heed wait!!!"));
          write(output, write_line91.all);
          deallocate (write_line91);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_clock_9_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_0_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal nios2_clock_9_in_endofpacket : IN STD_LOGIC;
                 signal nios2_clock_9_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_9_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_byteenable_nios2_clock_9_in : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_0_data_master_granted_nios2_clock_9_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_nios2_clock_9_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_nios2_clock_9_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_nios2_clock_9_in : OUT STD_LOGIC;
                 signal d1_nios2_clock_9_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_9_in_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_9_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_9_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_9_in_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal nios2_clock_9_in_read : OUT STD_LOGIC;
                 signal nios2_clock_9_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_9_in_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_9_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_clock_9_in_write : OUT STD_LOGIC;
                 signal nios2_clock_9_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity nios2_clock_9_in_arbitrator;


architecture europa of nios2_clock_9_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_byteenable_nios2_clock_9_in_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_data_master_byteenable_nios2_clock_9_in_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_nios2_clock_9_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_clock_9_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_byteenable_nios2_clock_9_in :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_0_data_master_granted_nios2_clock_9_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_nios2_clock_9_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_nios2_clock_9_in :  STD_LOGIC;
                signal internal_nios2_clock_9_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_9_in_allgrants :  STD_LOGIC;
                signal nios2_clock_9_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_clock_9_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_clock_9_in_any_continuerequest :  STD_LOGIC;
                signal nios2_clock_9_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_clock_9_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_9_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_9_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_9_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_clock_9_in_begins_xfer :  STD_LOGIC;
                signal nios2_clock_9_in_end_xfer :  STD_LOGIC;
                signal nios2_clock_9_in_firsttransfer :  STD_LOGIC;
                signal nios2_clock_9_in_grant_vector :  STD_LOGIC;
                signal nios2_clock_9_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_clock_9_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_clock_9_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_clock_9_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_clock_9_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_9_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_clock_9_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_clock_9_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_clock_9_in_waits_for_read :  STD_LOGIC;
                signal nios2_clock_9_in_waits_for_write :  STD_LOGIC;
                signal wait_for_nios2_clock_9_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_clock_9_in_end_xfer;
    end if;

  end process;

  nios2_clock_9_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_nios2_clock_9_in);
  --assign nios2_clock_9_in_readdata_from_sa = nios2_clock_9_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_9_in_readdata_from_sa <= nios2_clock_9_in_readdata;
  internal_cpu_0_data_master_requests_nios2_clock_9_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(24 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("0100000000000000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign nios2_clock_9_in_waitrequest_from_sa = nios2_clock_9_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_clock_9_in_waitrequest_from_sa <= nios2_clock_9_in_waitrequest;
  --nios2_clock_9_in_arb_share_counter set values, which is an e_mux
  nios2_clock_9_in_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_9_in)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001")), 2);
  --nios2_clock_9_in_non_bursting_master_requests mux, which is an e_mux
  nios2_clock_9_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_nios2_clock_9_in;
  --nios2_clock_9_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_clock_9_in_any_bursting_master_saved_grant <= std_logic'('0');
  --nios2_clock_9_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_clock_9_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_clock_9_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_9_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_clock_9_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_clock_9_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --nios2_clock_9_in_allgrants all slave grants, which is an e_mux
  nios2_clock_9_in_allgrants <= nios2_clock_9_in_grant_vector;
  --nios2_clock_9_in_end_xfer assignment, which is an e_assign
  nios2_clock_9_in_end_xfer <= NOT ((nios2_clock_9_in_waits_for_read OR nios2_clock_9_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_clock_9_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_clock_9_in <= nios2_clock_9_in_end_xfer AND (((NOT nios2_clock_9_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_clock_9_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_clock_9_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_clock_9_in AND nios2_clock_9_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_clock_9_in AND NOT nios2_clock_9_in_non_bursting_master_requests));
  --nios2_clock_9_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_9_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_9_in_arb_counter_enable) = '1' then 
        nios2_clock_9_in_arb_share_counter <= nios2_clock_9_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_9_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_9_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_clock_9_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_clock_9_in)) OR ((end_xfer_arb_share_counter_term_nios2_clock_9_in AND NOT nios2_clock_9_in_non_bursting_master_requests)))) = '1' then 
        nios2_clock_9_in_slavearbiterlockenable <= or_reduce(nios2_clock_9_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_0/data_master nios2_clock_9/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= nios2_clock_9_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --nios2_clock_9_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_clock_9_in_slavearbiterlockenable2 <= or_reduce(nios2_clock_9_in_arb_share_counter_next_value);
  --cpu_0/data_master nios2_clock_9/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= nios2_clock_9_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --nios2_clock_9_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_clock_9_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_nios2_clock_9_in <= internal_cpu_0_data_master_requests_nios2_clock_9_in AND NOT ((((cpu_0_data_master_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR (((NOT(or_reduce(internal_cpu_0_data_master_byteenable_nios2_clock_9_in))) AND cpu_0_data_master_write))));
  --local readdatavalid cpu_0_data_master_read_data_valid_nios2_clock_9_in, which is an e_mux
  cpu_0_data_master_read_data_valid_nios2_clock_9_in <= (internal_cpu_0_data_master_granted_nios2_clock_9_in AND cpu_0_data_master_read) AND NOT nios2_clock_9_in_waits_for_read;
  --nios2_clock_9_in_writedata mux, which is an e_mux
  nios2_clock_9_in_writedata <= cpu_0_data_master_dbs_write_16;
  --assign nios2_clock_9_in_endofpacket_from_sa = nios2_clock_9_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_clock_9_in_endofpacket_from_sa <= nios2_clock_9_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_nios2_clock_9_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_9_in;
  --cpu_0/data_master saved-grant nios2_clock_9/in, which is an e_assign
  cpu_0_data_master_saved_grant_nios2_clock_9_in <= internal_cpu_0_data_master_requests_nios2_clock_9_in;
  --allow new arb cycle for nios2_clock_9/in, which is an e_assign
  nios2_clock_9_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_clock_9_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_clock_9_in_master_qreq_vector <= std_logic'('1');
  --nios2_clock_9_in_reset_n assignment, which is an e_assign
  nios2_clock_9_in_reset_n <= reset_n;
  --nios2_clock_9_in_firsttransfer first transaction, which is an e_assign
  nios2_clock_9_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_clock_9_in_begins_xfer) = '1'), nios2_clock_9_in_unreg_firsttransfer, nios2_clock_9_in_reg_firsttransfer);
  --nios2_clock_9_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_clock_9_in_unreg_firsttransfer <= NOT ((nios2_clock_9_in_slavearbiterlockenable AND nios2_clock_9_in_any_continuerequest));
  --nios2_clock_9_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_9_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_clock_9_in_begins_xfer) = '1' then 
        nios2_clock_9_in_reg_firsttransfer <= nios2_clock_9_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_clock_9_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_clock_9_in_beginbursttransfer_internal <= nios2_clock_9_in_begins_xfer;
  --nios2_clock_9_in_read assignment, which is an e_mux
  nios2_clock_9_in_read <= internal_cpu_0_data_master_granted_nios2_clock_9_in AND cpu_0_data_master_read;
  --nios2_clock_9_in_write assignment, which is an e_mux
  nios2_clock_9_in_write <= internal_cpu_0_data_master_granted_nios2_clock_9_in AND cpu_0_data_master_write;
  --nios2_clock_9_in_address mux, which is an e_mux
  nios2_clock_9_in_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_0_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 23);
  --slaveid nios2_clock_9_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_clock_9_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 22);
  --d1_nios2_clock_9_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_clock_9_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_clock_9_in_end_xfer <= nios2_clock_9_in_end_xfer;
    end if;

  end process;

  --nios2_clock_9_in_waits_for_read in a cycle, which is an e_mux
  nios2_clock_9_in_waits_for_read <= nios2_clock_9_in_in_a_read_cycle AND internal_nios2_clock_9_in_waitrequest_from_sa;
  --nios2_clock_9_in_in_a_read_cycle assignment, which is an e_assign
  nios2_clock_9_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_nios2_clock_9_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_clock_9_in_in_a_read_cycle;
  --nios2_clock_9_in_waits_for_write in a cycle, which is an e_mux
  nios2_clock_9_in_waits_for_write <= nios2_clock_9_in_in_a_write_cycle AND internal_nios2_clock_9_in_waitrequest_from_sa;
  --nios2_clock_9_in_in_a_write_cycle assignment, which is an e_assign
  nios2_clock_9_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_nios2_clock_9_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_clock_9_in_in_a_write_cycle;
  wait_for_nios2_clock_9_in_counter <= std_logic'('0');
  --nios2_clock_9_in_byteenable byte enable port mux, which is an e_mux
  nios2_clock_9_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_nios2_clock_9_in)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_cpu_0_data_master_byteenable_nios2_clock_9_in)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  (cpu_0_data_master_byteenable_nios2_clock_9_in_segment_1(1), cpu_0_data_master_byteenable_nios2_clock_9_in_segment_1(0), cpu_0_data_master_byteenable_nios2_clock_9_in_segment_0(1), cpu_0_data_master_byteenable_nios2_clock_9_in_segment_0(0)) <= cpu_0_data_master_byteenable;
  internal_cpu_0_data_master_byteenable_nios2_clock_9_in <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_0_data_master_byteenable_nios2_clock_9_in_segment_0, cpu_0_data_master_byteenable_nios2_clock_9_in_segment_1);
  --vhdl renameroo for output signals
  cpu_0_data_master_byteenable_nios2_clock_9_in <= internal_cpu_0_data_master_byteenable_nios2_clock_9_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_nios2_clock_9_in <= internal_cpu_0_data_master_granted_nios2_clock_9_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_nios2_clock_9_in <= internal_cpu_0_data_master_qualified_request_nios2_clock_9_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_nios2_clock_9_in <= internal_cpu_0_data_master_requests_nios2_clock_9_in;
  --vhdl renameroo for output signals
  nios2_clock_9_in_waitrequest_from_sa <= internal_nios2_clock_9_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_clock_9/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_clock_9_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_clock_9_out_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_9_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_9_out_granted_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_9_out_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_9_out_read : IN STD_LOGIC;
                 signal nios2_clock_9_out_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal nios2_clock_9_out_requests_sdram_0_s1 : IN STD_LOGIC;
                 signal nios2_clock_9_out_write : IN STD_LOGIC;
                 signal nios2_clock_9_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_clock_9_out_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_9_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_9_out_reset_n : OUT STD_LOGIC;
                 signal nios2_clock_9_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_clock_9_out_arbitrator;


architecture europa of nios2_clock_9_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_clock_9_out_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal internal_nios2_clock_9_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_9_out_address_last_time :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_9_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_9_out_read_last_time :  STD_LOGIC;
                signal nios2_clock_9_out_run :  STD_LOGIC;
                signal nios2_clock_9_out_write_last_time :  STD_LOGIC;
                signal nios2_clock_9_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal r_3 :  STD_LOGIC;

begin

  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((nios2_clock_9_out_qualified_request_sdram_0_s1 OR nios2_clock_9_out_read_data_valid_sdram_0_s1) OR NOT nios2_clock_9_out_requests_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_9_out_granted_sdram_0_s1 OR NOT nios2_clock_9_out_qualified_request_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT nios2_clock_9_out_qualified_request_sdram_0_s1 OR NOT nios2_clock_9_out_read) OR ((nios2_clock_9_out_read_data_valid_sdram_0_s1 AND nios2_clock_9_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_clock_9_out_qualified_request_sdram_0_s1 OR NOT ((nios2_clock_9_out_read OR nios2_clock_9_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_0_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_9_out_read OR nios2_clock_9_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_clock_9_out_run <= r_3;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_clock_9_out_address_to_slave <= nios2_clock_9_out_address;
  --nios2_clock_9/out readdata mux, which is an e_mux
  nios2_clock_9_out_readdata <= sdram_0_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_clock_9_out_waitrequest <= NOT nios2_clock_9_out_run;
  --nios2_clock_9_out_reset_n assignment, which is an e_assign
  nios2_clock_9_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_clock_9_out_address_to_slave <= internal_nios2_clock_9_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_clock_9_out_waitrequest <= internal_nios2_clock_9_out_waitrequest;
--synthesis translate_off
    --nios2_clock_9_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_9_out_address_last_time <= std_logic_vector'("00000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_9_out_address_last_time <= nios2_clock_9_out_address;
      end if;

    end process;

    --nios2_clock_9/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_clock_9_out_waitrequest AND ((nios2_clock_9_out_read OR nios2_clock_9_out_write));
      end if;

    end process;

    --nios2_clock_9_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line92 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_9_out_address /= nios2_clock_9_out_address_last_time))))) = '1' then 
          write(write_line92, now);
          write(write_line92, string'(": "));
          write(write_line92, string'("nios2_clock_9_out_address did not heed wait!!!"));
          write(output, write_line92.all);
          deallocate (write_line92);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_9_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_9_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_clock_9_out_byteenable_last_time <= nios2_clock_9_out_byteenable;
      end if;

    end process;

    --nios2_clock_9_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line93 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_clock_9_out_byteenable /= nios2_clock_9_out_byteenable_last_time))))) = '1' then 
          write(write_line93, now);
          write(write_line93, string'(": "));
          write(write_line93, string'("nios2_clock_9_out_byteenable did not heed wait!!!"));
          write(output, write_line93.all);
          deallocate (write_line93);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_9_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_9_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_9_out_read_last_time <= nios2_clock_9_out_read;
      end if;

    end process;

    --nios2_clock_9_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line94 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_9_out_read) /= std_logic'(nios2_clock_9_out_read_last_time)))))) = '1' then 
          write(write_line94, now);
          write(write_line94, string'(": "));
          write(write_line94, string'("nios2_clock_9_out_read did not heed wait!!!"));
          write(output, write_line94.all);
          deallocate (write_line94);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_9_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_9_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_clock_9_out_write_last_time <= nios2_clock_9_out_write;
      end if;

    end process;

    --nios2_clock_9_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line95 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_clock_9_out_write) /= std_logic'(nios2_clock_9_out_write_last_time)))))) = '1' then 
          write(write_line95, now);
          write(write_line95, string'(": "));
          write(write_line95, string'("nios2_clock_9_out_write did not heed wait!!!"));
          write(output, write_line95.all);
          deallocate (write_line95);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_clock_9_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_clock_9_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_clock_9_out_writedata_last_time <= nios2_clock_9_out_writedata;
      end if;

    end process;

    --nios2_clock_9_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line96 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_clock_9_out_writedata /= nios2_clock_9_out_writedata_last_time)))) AND nios2_clock_9_out_write)) = '1' then 
          write(write_line96, now);
          write(write_line96, string'(": "));
          write(write_line96, string'("nios2_clock_9_out_writedata did not heed wait!!!"));
          write(output, write_line96.all);
          deallocate (write_line96);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity onchip_mem_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_0_out_read : IN STD_LOGIC;
                 signal nios2_clock_0_out_write : IN STD_LOGIC;
                 signal nios2_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_1_out_read : IN STD_LOGIC;
                 signal nios2_clock_1_out_write : IN STD_LOGIC;
                 signal nios2_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal onchip_mem_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_onchip_mem_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_0_out_granted_onchip_mem_s1 : OUT STD_LOGIC;
                 signal nios2_clock_0_out_qualified_request_onchip_mem_s1 : OUT STD_LOGIC;
                 signal nios2_clock_0_out_read_data_valid_onchip_mem_s1 : OUT STD_LOGIC;
                 signal nios2_clock_0_out_requests_onchip_mem_s1 : OUT STD_LOGIC;
                 signal nios2_clock_1_out_granted_onchip_mem_s1 : OUT STD_LOGIC;
                 signal nios2_clock_1_out_qualified_request_onchip_mem_s1 : OUT STD_LOGIC;
                 signal nios2_clock_1_out_read_data_valid_onchip_mem_s1 : OUT STD_LOGIC;
                 signal nios2_clock_1_out_requests_onchip_mem_s1 : OUT STD_LOGIC;
                 signal onchip_mem_s1_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal onchip_mem_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal onchip_mem_s1_chipselect : OUT STD_LOGIC;
                 signal onchip_mem_s1_clken : OUT STD_LOGIC;
                 signal onchip_mem_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal onchip_mem_s1_reset : OUT STD_LOGIC;
                 signal onchip_mem_s1_write : OUT STD_LOGIC;
                 signal onchip_mem_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity onchip_mem_s1_arbitrator;


architecture europa of onchip_mem_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_onchip_mem_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_0_out_granted_onchip_mem_s1 :  STD_LOGIC;
                signal internal_nios2_clock_0_out_qualified_request_onchip_mem_s1 :  STD_LOGIC;
                signal internal_nios2_clock_0_out_requests_onchip_mem_s1 :  STD_LOGIC;
                signal internal_nios2_clock_1_out_granted_onchip_mem_s1 :  STD_LOGIC;
                signal internal_nios2_clock_1_out_qualified_request_onchip_mem_s1 :  STD_LOGIC;
                signal internal_nios2_clock_1_out_requests_onchip_mem_s1 :  STD_LOGIC;
                signal last_cycle_nios2_clock_0_out_granted_slave_onchip_mem_s1 :  STD_LOGIC;
                signal last_cycle_nios2_clock_1_out_granted_slave_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_0_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_0_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_0_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register :  STD_LOGIC;
                signal nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register_in :  STD_LOGIC;
                signal nios2_clock_0_out_saved_grant_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_1_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_1_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_1_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register :  STD_LOGIC;
                signal nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register_in :  STD_LOGIC;
                signal nios2_clock_1_out_saved_grant_onchip_mem_s1 :  STD_LOGIC;
                signal onchip_mem_s1_allgrants :  STD_LOGIC;
                signal onchip_mem_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal onchip_mem_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal onchip_mem_s1_any_continuerequest :  STD_LOGIC;
                signal onchip_mem_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_mem_s1_arb_counter_enable :  STD_LOGIC;
                signal onchip_mem_s1_arb_share_counter :  STD_LOGIC;
                signal onchip_mem_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal onchip_mem_s1_arb_share_set_values :  STD_LOGIC;
                signal onchip_mem_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_mem_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal onchip_mem_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal onchip_mem_s1_begins_xfer :  STD_LOGIC;
                signal onchip_mem_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal onchip_mem_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_mem_s1_end_xfer :  STD_LOGIC;
                signal onchip_mem_s1_firsttransfer :  STD_LOGIC;
                signal onchip_mem_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_mem_s1_in_a_read_cycle :  STD_LOGIC;
                signal onchip_mem_s1_in_a_write_cycle :  STD_LOGIC;
                signal onchip_mem_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_mem_s1_non_bursting_master_requests :  STD_LOGIC;
                signal onchip_mem_s1_reg_firsttransfer :  STD_LOGIC;
                signal onchip_mem_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_mem_s1_slavearbiterlockenable :  STD_LOGIC;
                signal onchip_mem_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal onchip_mem_s1_unreg_firsttransfer :  STD_LOGIC;
                signal onchip_mem_s1_waits_for_read :  STD_LOGIC;
                signal onchip_mem_s1_waits_for_write :  STD_LOGIC;
                signal p1_nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register :  STD_LOGIC;
                signal p1_nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register :  STD_LOGIC;
                signal shifted_address_to_onchip_mem_s1_from_nios2_clock_0_out :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal shifted_address_to_onchip_mem_s1_from_nios2_clock_1_out :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal wait_for_onchip_mem_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT onchip_mem_s1_end_xfer;
    end if;

  end process;

  onchip_mem_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_nios2_clock_0_out_qualified_request_onchip_mem_s1 OR internal_nios2_clock_1_out_qualified_request_onchip_mem_s1));
  --assign onchip_mem_s1_readdata_from_sa = onchip_mem_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  onchip_mem_s1_readdata_from_sa <= onchip_mem_s1_readdata;
  internal_nios2_clock_0_out_requests_onchip_mem_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_0_out_read OR nios2_clock_0_out_write)))))));
  --onchip_mem_s1_arb_share_counter set values, which is an e_mux
  onchip_mem_s1_arb_share_set_values <= std_logic'('1');
  --onchip_mem_s1_non_bursting_master_requests mux, which is an e_mux
  onchip_mem_s1_non_bursting_master_requests <= ((internal_nios2_clock_0_out_requests_onchip_mem_s1 OR internal_nios2_clock_1_out_requests_onchip_mem_s1) OR internal_nios2_clock_0_out_requests_onchip_mem_s1) OR internal_nios2_clock_1_out_requests_onchip_mem_s1;
  --onchip_mem_s1_any_bursting_master_saved_grant mux, which is an e_mux
  onchip_mem_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --onchip_mem_s1_arb_share_counter_next_value assignment, which is an e_assign
  onchip_mem_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(onchip_mem_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_mem_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(onchip_mem_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_mem_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --onchip_mem_s1_allgrants all slave grants, which is an e_mux
  onchip_mem_s1_allgrants <= (((or_reduce(onchip_mem_s1_grant_vector)) OR (or_reduce(onchip_mem_s1_grant_vector))) OR (or_reduce(onchip_mem_s1_grant_vector))) OR (or_reduce(onchip_mem_s1_grant_vector));
  --onchip_mem_s1_end_xfer assignment, which is an e_assign
  onchip_mem_s1_end_xfer <= NOT ((onchip_mem_s1_waits_for_read OR onchip_mem_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_onchip_mem_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_onchip_mem_s1 <= onchip_mem_s1_end_xfer AND (((NOT onchip_mem_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --onchip_mem_s1_arb_share_counter arbitration counter enable, which is an e_assign
  onchip_mem_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_onchip_mem_s1 AND onchip_mem_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_onchip_mem_s1 AND NOT onchip_mem_s1_non_bursting_master_requests));
  --onchip_mem_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_mem_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_mem_s1_arb_counter_enable) = '1' then 
        onchip_mem_s1_arb_share_counter <= onchip_mem_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --onchip_mem_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_mem_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(onchip_mem_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_onchip_mem_s1)) OR ((end_xfer_arb_share_counter_term_onchip_mem_s1 AND NOT onchip_mem_s1_non_bursting_master_requests)))) = '1' then 
        onchip_mem_s1_slavearbiterlockenable <= onchip_mem_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_0/out onchip_mem/s1 arbiterlock, which is an e_assign
  nios2_clock_0_out_arbiterlock <= onchip_mem_s1_slavearbiterlockenable AND nios2_clock_0_out_continuerequest;
  --onchip_mem_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  onchip_mem_s1_slavearbiterlockenable2 <= onchip_mem_s1_arb_share_counter_next_value;
  --nios2_clock_0/out onchip_mem/s1 arbiterlock2, which is an e_assign
  nios2_clock_0_out_arbiterlock2 <= onchip_mem_s1_slavearbiterlockenable2 AND nios2_clock_0_out_continuerequest;
  --nios2_clock_1/out onchip_mem/s1 arbiterlock, which is an e_assign
  nios2_clock_1_out_arbiterlock <= onchip_mem_s1_slavearbiterlockenable AND nios2_clock_1_out_continuerequest;
  --nios2_clock_1/out onchip_mem/s1 arbiterlock2, which is an e_assign
  nios2_clock_1_out_arbiterlock2 <= onchip_mem_s1_slavearbiterlockenable2 AND nios2_clock_1_out_continuerequest;
  --nios2_clock_1/out granted onchip_mem/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_clock_1_out_granted_slave_onchip_mem_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_clock_1_out_granted_slave_onchip_mem_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_clock_1_out_saved_grant_onchip_mem_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((onchip_mem_s1_arbitration_holdoff_internal OR NOT internal_nios2_clock_1_out_requests_onchip_mem_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_clock_1_out_granted_slave_onchip_mem_s1))))));
    end if;

  end process;

  --nios2_clock_1_out_continuerequest continued request, which is an e_mux
  nios2_clock_1_out_continuerequest <= last_cycle_nios2_clock_1_out_granted_slave_onchip_mem_s1 AND internal_nios2_clock_1_out_requests_onchip_mem_s1;
  --onchip_mem_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  onchip_mem_s1_any_continuerequest <= nios2_clock_1_out_continuerequest OR nios2_clock_0_out_continuerequest;
  internal_nios2_clock_0_out_qualified_request_onchip_mem_s1 <= internal_nios2_clock_0_out_requests_onchip_mem_s1 AND NOT ((((nios2_clock_0_out_read AND (nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register))) OR nios2_clock_1_out_arbiterlock));
  --nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register_in <= ((internal_nios2_clock_0_out_granted_onchip_mem_s1 AND nios2_clock_0_out_read) AND NOT onchip_mem_s1_waits_for_read) AND NOT (nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register);
  --shift register p1 nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register) & A_ToStdLogicVector(nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register_in)));
  --nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register <= p1_nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register;
    end if;

  end process;

  --local readdatavalid nios2_clock_0_out_read_data_valid_onchip_mem_s1, which is an e_mux
  nios2_clock_0_out_read_data_valid_onchip_mem_s1 <= nios2_clock_0_out_read_data_valid_onchip_mem_s1_shift_register;
  --onchip_mem_s1_writedata mux, which is an e_mux
  onchip_mem_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_nios2_clock_0_out_granted_onchip_mem_s1)) = '1'), nios2_clock_0_out_writedata, nios2_clock_1_out_writedata);
  --mux onchip_mem_s1_clken, which is an e_mux
  onchip_mem_s1_clken <= std_logic'('1');
  internal_nios2_clock_1_out_requests_onchip_mem_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_1_out_read OR nios2_clock_1_out_write)))))));
  --nios2_clock_0/out granted onchip_mem/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_clock_0_out_granted_slave_onchip_mem_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_clock_0_out_granted_slave_onchip_mem_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_clock_0_out_saved_grant_onchip_mem_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((onchip_mem_s1_arbitration_holdoff_internal OR NOT internal_nios2_clock_0_out_requests_onchip_mem_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_clock_0_out_granted_slave_onchip_mem_s1))))));
    end if;

  end process;

  --nios2_clock_0_out_continuerequest continued request, which is an e_mux
  nios2_clock_0_out_continuerequest <= last_cycle_nios2_clock_0_out_granted_slave_onchip_mem_s1 AND internal_nios2_clock_0_out_requests_onchip_mem_s1;
  internal_nios2_clock_1_out_qualified_request_onchip_mem_s1 <= internal_nios2_clock_1_out_requests_onchip_mem_s1 AND NOT ((((nios2_clock_1_out_read AND (nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register))) OR nios2_clock_0_out_arbiterlock));
  --nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register_in <= ((internal_nios2_clock_1_out_granted_onchip_mem_s1 AND nios2_clock_1_out_read) AND NOT onchip_mem_s1_waits_for_read) AND NOT (nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register);
  --shift register p1 nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register) & A_ToStdLogicVector(nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register_in)));
  --nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register <= p1_nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register;
    end if;

  end process;

  --local readdatavalid nios2_clock_1_out_read_data_valid_onchip_mem_s1, which is an e_mux
  nios2_clock_1_out_read_data_valid_onchip_mem_s1 <= nios2_clock_1_out_read_data_valid_onchip_mem_s1_shift_register;
  --allow new arb cycle for onchip_mem/s1, which is an e_assign
  onchip_mem_s1_allow_new_arb_cycle <= NOT nios2_clock_0_out_arbiterlock AND NOT nios2_clock_1_out_arbiterlock;
  --nios2_clock_1/out assignment into master qualified-requests vector for onchip_mem/s1, which is an e_assign
  onchip_mem_s1_master_qreq_vector(0) <= internal_nios2_clock_1_out_qualified_request_onchip_mem_s1;
  --nios2_clock_1/out grant onchip_mem/s1, which is an e_assign
  internal_nios2_clock_1_out_granted_onchip_mem_s1 <= onchip_mem_s1_grant_vector(0);
  --nios2_clock_1/out saved-grant onchip_mem/s1, which is an e_assign
  nios2_clock_1_out_saved_grant_onchip_mem_s1 <= onchip_mem_s1_arb_winner(0) AND internal_nios2_clock_1_out_requests_onchip_mem_s1;
  --nios2_clock_0/out assignment into master qualified-requests vector for onchip_mem/s1, which is an e_assign
  onchip_mem_s1_master_qreq_vector(1) <= internal_nios2_clock_0_out_qualified_request_onchip_mem_s1;
  --nios2_clock_0/out grant onchip_mem/s1, which is an e_assign
  internal_nios2_clock_0_out_granted_onchip_mem_s1 <= onchip_mem_s1_grant_vector(1);
  --nios2_clock_0/out saved-grant onchip_mem/s1, which is an e_assign
  nios2_clock_0_out_saved_grant_onchip_mem_s1 <= onchip_mem_s1_arb_winner(1) AND internal_nios2_clock_0_out_requests_onchip_mem_s1;
  --onchip_mem/s1 chosen-master double-vector, which is an e_assign
  onchip_mem_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((onchip_mem_s1_master_qreq_vector & onchip_mem_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT onchip_mem_s1_master_qreq_vector & NOT onchip_mem_s1_master_qreq_vector))) + (std_logic_vector'("000") & (onchip_mem_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  onchip_mem_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((onchip_mem_s1_allow_new_arb_cycle AND or_reduce(onchip_mem_s1_grant_vector)))) = '1'), onchip_mem_s1_grant_vector, onchip_mem_s1_saved_chosen_master_vector);
  --saved onchip_mem_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_mem_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_mem_s1_allow_new_arb_cycle) = '1' then 
        onchip_mem_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(onchip_mem_s1_grant_vector)) = '1'), onchip_mem_s1_grant_vector, onchip_mem_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  onchip_mem_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((onchip_mem_s1_chosen_master_double_vector(1) OR onchip_mem_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((onchip_mem_s1_chosen_master_double_vector(0) OR onchip_mem_s1_chosen_master_double_vector(2)))));
  --onchip_mem/s1 chosen master rotated left, which is an e_assign
  onchip_mem_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(onchip_mem_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(onchip_mem_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --onchip_mem/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_mem_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(onchip_mem_s1_grant_vector)) = '1' then 
        onchip_mem_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(onchip_mem_s1_end_xfer) = '1'), onchip_mem_s1_chosen_master_rot_left, onchip_mem_s1_grant_vector);
      end if;
    end if;

  end process;

  --~onchip_mem_s1_reset assignment, which is an e_assign
  onchip_mem_s1_reset <= NOT reset_n;
  onchip_mem_s1_chipselect <= internal_nios2_clock_0_out_granted_onchip_mem_s1 OR internal_nios2_clock_1_out_granted_onchip_mem_s1;
  --onchip_mem_s1_firsttransfer first transaction, which is an e_assign
  onchip_mem_s1_firsttransfer <= A_WE_StdLogic((std_logic'(onchip_mem_s1_begins_xfer) = '1'), onchip_mem_s1_unreg_firsttransfer, onchip_mem_s1_reg_firsttransfer);
  --onchip_mem_s1_unreg_firsttransfer first transaction, which is an e_assign
  onchip_mem_s1_unreg_firsttransfer <= NOT ((onchip_mem_s1_slavearbiterlockenable AND onchip_mem_s1_any_continuerequest));
  --onchip_mem_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_mem_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_mem_s1_begins_xfer) = '1' then 
        onchip_mem_s1_reg_firsttransfer <= onchip_mem_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --onchip_mem_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  onchip_mem_s1_beginbursttransfer_internal <= onchip_mem_s1_begins_xfer;
  --onchip_mem_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  onchip_mem_s1_arbitration_holdoff_internal <= onchip_mem_s1_begins_xfer AND onchip_mem_s1_firsttransfer;
  --onchip_mem_s1_write assignment, which is an e_mux
  onchip_mem_s1_write <= ((internal_nios2_clock_0_out_granted_onchip_mem_s1 AND nios2_clock_0_out_write)) OR ((internal_nios2_clock_1_out_granted_onchip_mem_s1 AND nios2_clock_1_out_write));
  shifted_address_to_onchip_mem_s1_from_nios2_clock_0_out <= nios2_clock_0_out_address_to_slave;
  --onchip_mem_s1_address mux, which is an e_mux
  onchip_mem_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_clock_0_out_granted_onchip_mem_s1)) = '1'), (A_SRL(shifted_address_to_onchip_mem_s1_from_nios2_clock_0_out,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_onchip_mem_s1_from_nios2_clock_1_out,std_logic_vector'("00000000000000000000000000000010")))), 13);
  shifted_address_to_onchip_mem_s1_from_nios2_clock_1_out <= nios2_clock_1_out_address_to_slave;
  --d1_onchip_mem_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_onchip_mem_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_onchip_mem_s1_end_xfer <= onchip_mem_s1_end_xfer;
    end if;

  end process;

  --onchip_mem_s1_waits_for_read in a cycle, which is an e_mux
  onchip_mem_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_mem_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --onchip_mem_s1_in_a_read_cycle assignment, which is an e_assign
  onchip_mem_s1_in_a_read_cycle <= ((internal_nios2_clock_0_out_granted_onchip_mem_s1 AND nios2_clock_0_out_read)) OR ((internal_nios2_clock_1_out_granted_onchip_mem_s1 AND nios2_clock_1_out_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= onchip_mem_s1_in_a_read_cycle;
  --onchip_mem_s1_waits_for_write in a cycle, which is an e_mux
  onchip_mem_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_mem_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --onchip_mem_s1_in_a_write_cycle assignment, which is an e_assign
  onchip_mem_s1_in_a_write_cycle <= ((internal_nios2_clock_0_out_granted_onchip_mem_s1 AND nios2_clock_0_out_write)) OR ((internal_nios2_clock_1_out_granted_onchip_mem_s1 AND nios2_clock_1_out_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= onchip_mem_s1_in_a_write_cycle;
  wait_for_onchip_mem_s1_counter <= std_logic'('0');
  --onchip_mem_s1_byteenable byte enable port mux, which is an e_mux
  onchip_mem_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_clock_0_out_granted_onchip_mem_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_clock_0_out_byteenable)), A_WE_StdLogicVector((std_logic'((internal_nios2_clock_1_out_granted_onchip_mem_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_clock_1_out_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --vhdl renameroo for output signals
  nios2_clock_0_out_granted_onchip_mem_s1 <= internal_nios2_clock_0_out_granted_onchip_mem_s1;
  --vhdl renameroo for output signals
  nios2_clock_0_out_qualified_request_onchip_mem_s1 <= internal_nios2_clock_0_out_qualified_request_onchip_mem_s1;
  --vhdl renameroo for output signals
  nios2_clock_0_out_requests_onchip_mem_s1 <= internal_nios2_clock_0_out_requests_onchip_mem_s1;
  --vhdl renameroo for output signals
  nios2_clock_1_out_granted_onchip_mem_s1 <= internal_nios2_clock_1_out_granted_onchip_mem_s1;
  --vhdl renameroo for output signals
  nios2_clock_1_out_qualified_request_onchip_mem_s1 <= internal_nios2_clock_1_out_qualified_request_onchip_mem_s1;
  --vhdl renameroo for output signals
  nios2_clock_1_out_requests_onchip_mem_s1 <= internal_nios2_clock_1_out_requests_onchip_mem_s1;
--synthesis translate_off
    --onchip_mem/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line97 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_clock_0_out_granted_onchip_mem_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_clock_1_out_granted_onchip_mem_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line97, now);
          write(write_line97, string'(": "));
          write(write_line97, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line97.all);
          deallocate (write_line97);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line98 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_clock_0_out_saved_grant_onchip_mem_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_clock_1_out_saved_grant_onchip_mem_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line98, now);
          write(write_line98, string'(": "));
          write(write_line98, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line98.all);
          deallocate (write_line98);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sample_and_hold_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_17_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_17_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_17_out_read : IN STD_LOGIC;
                 signal nios2_clock_17_out_write : IN STD_LOGIC;
                 signal nios2_clock_17_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sample_and_hold_pio_s1_readdata : IN STD_LOGIC;

              -- outputs:
                 signal d1_sample_and_hold_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_17_out_granted_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_17_out_requests_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                 signal sample_and_hold_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sample_and_hold_pio_s1_chipselect : OUT STD_LOGIC;
                 signal sample_and_hold_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal sample_and_hold_pio_s1_reset_n : OUT STD_LOGIC;
                 signal sample_and_hold_pio_s1_write_n : OUT STD_LOGIC;
                 signal sample_and_hold_pio_s1_writedata : OUT STD_LOGIC
              );
end entity sample_and_hold_pio_s1_arbitrator;


architecture europa of sample_and_hold_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_17_out_granted_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_17_out_requests_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal nios2_clock_17_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_17_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_17_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_17_out_saved_grant_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal sample_and_hold_pio_s1_allgrants :  STD_LOGIC;
                signal sample_and_hold_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sample_and_hold_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sample_and_hold_pio_s1_any_continuerequest :  STD_LOGIC;
                signal sample_and_hold_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal sample_and_hold_pio_s1_arb_share_counter :  STD_LOGIC;
                signal sample_and_hold_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sample_and_hold_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal sample_and_hold_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sample_and_hold_pio_s1_begins_xfer :  STD_LOGIC;
                signal sample_and_hold_pio_s1_end_xfer :  STD_LOGIC;
                signal sample_and_hold_pio_s1_firsttransfer :  STD_LOGIC;
                signal sample_and_hold_pio_s1_grant_vector :  STD_LOGIC;
                signal sample_and_hold_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal sample_and_hold_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal sample_and_hold_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal sample_and_hold_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sample_and_hold_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal sample_and_hold_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sample_and_hold_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sample_and_hold_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sample_and_hold_pio_s1_waits_for_read :  STD_LOGIC;
                signal sample_and_hold_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sample_and_hold_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sample_and_hold_pio_s1_end_xfer;
    end if;

  end process;

  sample_and_hold_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1);
  --assign sample_and_hold_pio_s1_readdata_from_sa = sample_and_hold_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sample_and_hold_pio_s1_readdata_from_sa <= sample_and_hold_pio_s1_readdata;
  internal_nios2_clock_17_out_requests_sample_and_hold_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_17_out_read OR nios2_clock_17_out_write)))))));
  --sample_and_hold_pio_s1_arb_share_counter set values, which is an e_mux
  sample_and_hold_pio_s1_arb_share_set_values <= std_logic'('1');
  --sample_and_hold_pio_s1_non_bursting_master_requests mux, which is an e_mux
  sample_and_hold_pio_s1_non_bursting_master_requests <= internal_nios2_clock_17_out_requests_sample_and_hold_pio_s1;
  --sample_and_hold_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sample_and_hold_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sample_and_hold_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  sample_and_hold_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sample_and_hold_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sample_and_hold_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sample_and_hold_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sample_and_hold_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sample_and_hold_pio_s1_allgrants all slave grants, which is an e_mux
  sample_and_hold_pio_s1_allgrants <= sample_and_hold_pio_s1_grant_vector;
  --sample_and_hold_pio_s1_end_xfer assignment, which is an e_assign
  sample_and_hold_pio_s1_end_xfer <= NOT ((sample_and_hold_pio_s1_waits_for_read OR sample_and_hold_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sample_and_hold_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sample_and_hold_pio_s1 <= sample_and_hold_pio_s1_end_xfer AND (((NOT sample_and_hold_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sample_and_hold_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sample_and_hold_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sample_and_hold_pio_s1 AND sample_and_hold_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sample_and_hold_pio_s1 AND NOT sample_and_hold_pio_s1_non_bursting_master_requests));
  --sample_and_hold_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sample_and_hold_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sample_and_hold_pio_s1_arb_counter_enable) = '1' then 
        sample_and_hold_pio_s1_arb_share_counter <= sample_and_hold_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sample_and_hold_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sample_and_hold_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sample_and_hold_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sample_and_hold_pio_s1)) OR ((end_xfer_arb_share_counter_term_sample_and_hold_pio_s1 AND NOT sample_and_hold_pio_s1_non_bursting_master_requests)))) = '1' then 
        sample_and_hold_pio_s1_slavearbiterlockenable <= sample_and_hold_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_17/out sample_and_hold_pio/s1 arbiterlock, which is an e_assign
  nios2_clock_17_out_arbiterlock <= sample_and_hold_pio_s1_slavearbiterlockenable AND nios2_clock_17_out_continuerequest;
  --sample_and_hold_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sample_and_hold_pio_s1_slavearbiterlockenable2 <= sample_and_hold_pio_s1_arb_share_counter_next_value;
  --nios2_clock_17/out sample_and_hold_pio/s1 arbiterlock2, which is an e_assign
  nios2_clock_17_out_arbiterlock2 <= sample_and_hold_pio_s1_slavearbiterlockenable2 AND nios2_clock_17_out_continuerequest;
  --sample_and_hold_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sample_and_hold_pio_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_17_out_continuerequest continued request, which is an e_assign
  nios2_clock_17_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 <= internal_nios2_clock_17_out_requests_sample_and_hold_pio_s1;
  --sample_and_hold_pio_s1_writedata mux, which is an e_mux
  sample_and_hold_pio_s1_writedata <= nios2_clock_17_out_writedata(0);
  --master is always granted when requested
  internal_nios2_clock_17_out_granted_sample_and_hold_pio_s1 <= internal_nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1;
  --nios2_clock_17/out saved-grant sample_and_hold_pio/s1, which is an e_assign
  nios2_clock_17_out_saved_grant_sample_and_hold_pio_s1 <= internal_nios2_clock_17_out_requests_sample_and_hold_pio_s1;
  --allow new arb cycle for sample_and_hold_pio/s1, which is an e_assign
  sample_and_hold_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sample_and_hold_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sample_and_hold_pio_s1_master_qreq_vector <= std_logic'('1');
  --sample_and_hold_pio_s1_reset_n assignment, which is an e_assign
  sample_and_hold_pio_s1_reset_n <= reset_n;
  sample_and_hold_pio_s1_chipselect <= internal_nios2_clock_17_out_granted_sample_and_hold_pio_s1;
  --sample_and_hold_pio_s1_firsttransfer first transaction, which is an e_assign
  sample_and_hold_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sample_and_hold_pio_s1_begins_xfer) = '1'), sample_and_hold_pio_s1_unreg_firsttransfer, sample_and_hold_pio_s1_reg_firsttransfer);
  --sample_and_hold_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  sample_and_hold_pio_s1_unreg_firsttransfer <= NOT ((sample_and_hold_pio_s1_slavearbiterlockenable AND sample_and_hold_pio_s1_any_continuerequest));
  --sample_and_hold_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sample_and_hold_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sample_and_hold_pio_s1_begins_xfer) = '1' then 
        sample_and_hold_pio_s1_reg_firsttransfer <= sample_and_hold_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sample_and_hold_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sample_and_hold_pio_s1_beginbursttransfer_internal <= sample_and_hold_pio_s1_begins_xfer;
  --~sample_and_hold_pio_s1_write_n assignment, which is an e_mux
  sample_and_hold_pio_s1_write_n <= NOT ((internal_nios2_clock_17_out_granted_sample_and_hold_pio_s1 AND nios2_clock_17_out_write));
  --sample_and_hold_pio_s1_address mux, which is an e_mux
  sample_and_hold_pio_s1_address <= nios2_clock_17_out_nativeaddress;
  --d1_sample_and_hold_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sample_and_hold_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sample_and_hold_pio_s1_end_xfer <= sample_and_hold_pio_s1_end_xfer;
    end if;

  end process;

  --sample_and_hold_pio_s1_waits_for_read in a cycle, which is an e_mux
  sample_and_hold_pio_s1_waits_for_read <= sample_and_hold_pio_s1_in_a_read_cycle AND sample_and_hold_pio_s1_begins_xfer;
  --sample_and_hold_pio_s1_in_a_read_cycle assignment, which is an e_assign
  sample_and_hold_pio_s1_in_a_read_cycle <= internal_nios2_clock_17_out_granted_sample_and_hold_pio_s1 AND nios2_clock_17_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sample_and_hold_pio_s1_in_a_read_cycle;
  --sample_and_hold_pio_s1_waits_for_write in a cycle, which is an e_mux
  sample_and_hold_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sample_and_hold_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sample_and_hold_pio_s1_in_a_write_cycle assignment, which is an e_assign
  sample_and_hold_pio_s1_in_a_write_cycle <= internal_nios2_clock_17_out_granted_sample_and_hold_pio_s1 AND nios2_clock_17_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sample_and_hold_pio_s1_in_a_write_cycle;
  wait_for_sample_and_hold_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_17_out_granted_sample_and_hold_pio_s1 <= internal_nios2_clock_17_out_granted_sample_and_hold_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 <= internal_nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_17_out_requests_sample_and_hold_pio_s1 <= internal_nios2_clock_17_out_requests_sample_and_hold_pio_s1;
--synthesis translate_off
    --sample_and_hold_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1_module;


architecture europa of rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_5;
  empty <= NOT(full_0);
  full_6 <= std_logic'('0');
  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1_module;


architecture europa of rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_5;
  empty <= NOT(full_0);
  full_6 <= std_logic'('0');
  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sdram_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_8_out_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_8_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_8_out_read : IN STD_LOGIC;
                 signal nios2_clock_8_out_write : IN STD_LOGIC;
                 signal nios2_clock_8_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_clock_9_out_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal nios2_clock_9_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_9_out_read : IN STD_LOGIC;
                 signal nios2_clock_9_out_write : IN STD_LOGIC;
                 signal nios2_clock_9_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_0_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_0_s1_readdatavalid : IN STD_LOGIC;
                 signal sdram_0_s1_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal d1_sdram_0_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_8_out_granted_sdram_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_8_out_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_8_out_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                 signal nios2_clock_8_out_requests_sdram_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_9_out_granted_sdram_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_9_out_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_9_out_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                 signal nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                 signal nios2_clock_9_out_requests_sdram_0_s1 : OUT STD_LOGIC;
                 signal sdram_0_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal sdram_0_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sdram_0_s1_chipselect : OUT STD_LOGIC;
                 signal sdram_0_s1_read_n : OUT STD_LOGIC;
                 signal sdram_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_0_s1_reset_n : OUT STD_LOGIC;
                 signal sdram_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal sdram_0_s1_write_n : OUT STD_LOGIC;
                 signal sdram_0_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sdram_0_s1_arbitrator;


architecture europa of sdram_0_s1_arbitrator is
component rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1_module;

component rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sdram_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_8_out_granted_sdram_0_s1 :  STD_LOGIC;
                signal internal_nios2_clock_8_out_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal internal_nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register :  STD_LOGIC;
                signal internal_nios2_clock_8_out_requests_sdram_0_s1 :  STD_LOGIC;
                signal internal_nios2_clock_9_out_granted_sdram_0_s1 :  STD_LOGIC;
                signal internal_nios2_clock_9_out_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal internal_nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register :  STD_LOGIC;
                signal internal_nios2_clock_9_out_requests_sdram_0_s1 :  STD_LOGIC;
                signal internal_sdram_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_nios2_clock_8_out_granted_slave_sdram_0_s1 :  STD_LOGIC;
                signal last_cycle_nios2_clock_9_out_granted_slave_sdram_0_s1 :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal nios2_clock_8_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_8_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_8_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_8_out_rdv_fifo_empty_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_8_out_rdv_fifo_output_from_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_8_out_saved_grant_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_9_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_9_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_9_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_9_out_rdv_fifo_empty_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_9_out_rdv_fifo_output_from_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_9_out_saved_grant_sdram_0_s1 :  STD_LOGIC;
                signal sdram_0_s1_allgrants :  STD_LOGIC;
                signal sdram_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sdram_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sdram_0_s1_any_continuerequest :  STD_LOGIC;
                signal sdram_0_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_arb_counter_enable :  STD_LOGIC;
                signal sdram_0_s1_arb_share_counter :  STD_LOGIC;
                signal sdram_0_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sdram_0_s1_arb_share_set_values :  STD_LOGIC;
                signal sdram_0_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal sdram_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sdram_0_s1_begins_xfer :  STD_LOGIC;
                signal sdram_0_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_0_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_end_xfer :  STD_LOGIC;
                signal sdram_0_s1_firsttransfer :  STD_LOGIC;
                signal sdram_0_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal sdram_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal sdram_0_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal sdram_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sdram_0_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal sdram_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal sdram_0_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sdram_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sdram_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sdram_0_s1_waits_for_read :  STD_LOGIC;
                signal sdram_0_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sdram_0_s1_from_nios2_clock_8_out :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal shifted_address_to_sdram_0_s1_from_nios2_clock_9_out :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal wait_for_sdram_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sdram_0_s1_end_xfer;
    end if;

  end process;

  sdram_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_nios2_clock_8_out_qualified_request_sdram_0_s1 OR internal_nios2_clock_9_out_qualified_request_sdram_0_s1));
  --assign sdram_0_s1_readdata_from_sa = sdram_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_0_s1_readdata_from_sa <= sdram_0_s1_readdata;
  internal_nios2_clock_8_out_requests_sdram_0_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_8_out_read OR nios2_clock_8_out_write)))))));
  --assign sdram_0_s1_waitrequest_from_sa = sdram_0_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_sdram_0_s1_waitrequest_from_sa <= sdram_0_s1_waitrequest;
  --assign sdram_0_s1_readdatavalid_from_sa = sdram_0_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_0_s1_readdatavalid_from_sa <= sdram_0_s1_readdatavalid;
  --sdram_0_s1_arb_share_counter set values, which is an e_mux
  sdram_0_s1_arb_share_set_values <= std_logic'('1');
  --sdram_0_s1_non_bursting_master_requests mux, which is an e_mux
  sdram_0_s1_non_bursting_master_requests <= ((internal_nios2_clock_8_out_requests_sdram_0_s1 OR internal_nios2_clock_9_out_requests_sdram_0_s1) OR internal_nios2_clock_8_out_requests_sdram_0_s1) OR internal_nios2_clock_9_out_requests_sdram_0_s1;
  --sdram_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sdram_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sdram_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  sdram_0_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sdram_0_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_0_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sdram_0_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_0_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sdram_0_s1_allgrants all slave grants, which is an e_mux
  sdram_0_s1_allgrants <= (((or_reduce(sdram_0_s1_grant_vector)) OR (or_reduce(sdram_0_s1_grant_vector))) OR (or_reduce(sdram_0_s1_grant_vector))) OR (or_reduce(sdram_0_s1_grant_vector));
  --sdram_0_s1_end_xfer assignment, which is an e_assign
  sdram_0_s1_end_xfer <= NOT ((sdram_0_s1_waits_for_read OR sdram_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sdram_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sdram_0_s1 <= sdram_0_s1_end_xfer AND (((NOT sdram_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sdram_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sdram_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sdram_0_s1 AND sdram_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sdram_0_s1 AND NOT sdram_0_s1_non_bursting_master_requests));
  --sdram_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_0_s1_arb_counter_enable) = '1' then 
        sdram_0_s1_arb_share_counter <= sdram_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sdram_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sdram_0_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_sdram_0_s1)) OR ((end_xfer_arb_share_counter_term_sdram_0_s1 AND NOT sdram_0_s1_non_bursting_master_requests)))) = '1' then 
        sdram_0_s1_slavearbiterlockenable <= sdram_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_8/out sdram_0/s1 arbiterlock, which is an e_assign
  nios2_clock_8_out_arbiterlock <= sdram_0_s1_slavearbiterlockenable AND nios2_clock_8_out_continuerequest;
  --sdram_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sdram_0_s1_slavearbiterlockenable2 <= sdram_0_s1_arb_share_counter_next_value;
  --nios2_clock_8/out sdram_0/s1 arbiterlock2, which is an e_assign
  nios2_clock_8_out_arbiterlock2 <= sdram_0_s1_slavearbiterlockenable2 AND nios2_clock_8_out_continuerequest;
  --nios2_clock_9/out sdram_0/s1 arbiterlock, which is an e_assign
  nios2_clock_9_out_arbiterlock <= sdram_0_s1_slavearbiterlockenable AND nios2_clock_9_out_continuerequest;
  --nios2_clock_9/out sdram_0/s1 arbiterlock2, which is an e_assign
  nios2_clock_9_out_arbiterlock2 <= sdram_0_s1_slavearbiterlockenable2 AND nios2_clock_9_out_continuerequest;
  --nios2_clock_9/out granted sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_clock_9_out_granted_slave_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_clock_9_out_granted_slave_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_clock_9_out_saved_grant_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_0_s1_arbitration_holdoff_internal OR NOT internal_nios2_clock_9_out_requests_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_clock_9_out_granted_slave_sdram_0_s1))))));
    end if;

  end process;

  --nios2_clock_9_out_continuerequest continued request, which is an e_mux
  nios2_clock_9_out_continuerequest <= last_cycle_nios2_clock_9_out_granted_slave_sdram_0_s1 AND internal_nios2_clock_9_out_requests_sdram_0_s1;
  --sdram_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  sdram_0_s1_any_continuerequest <= nios2_clock_9_out_continuerequest OR nios2_clock_8_out_continuerequest;
  internal_nios2_clock_8_out_qualified_request_sdram_0_s1 <= internal_nios2_clock_8_out_requests_sdram_0_s1 AND NOT ((((nios2_clock_8_out_read AND (internal_nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register))) OR nios2_clock_9_out_arbiterlock));
  --unique name for sdram_0_s1_move_on_to_next_transaction, which is an e_assign
  sdram_0_s1_move_on_to_next_transaction <= sdram_0_s1_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1 : rdv_fifo_for_nios2_clock_8_out_to_sdram_0_s1_module
    port map(
      data_out => nios2_clock_8_out_rdv_fifo_output_from_sdram_0_s1,
      empty => open,
      fifo_contains_ones_n => nios2_clock_8_out_rdv_fifo_empty_sdram_0_s1,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => internal_nios2_clock_8_out_granted_sdram_0_s1,
      read => sdram_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= in_a_read_cycle AND NOT sdram_0_s1_waits_for_read;

  internal_nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register <= NOT nios2_clock_8_out_rdv_fifo_empty_sdram_0_s1;
  --local readdatavalid nios2_clock_8_out_read_data_valid_sdram_0_s1, which is an e_mux
  nios2_clock_8_out_read_data_valid_sdram_0_s1 <= ((sdram_0_s1_readdatavalid_from_sa AND nios2_clock_8_out_rdv_fifo_output_from_sdram_0_s1)) AND NOT nios2_clock_8_out_rdv_fifo_empty_sdram_0_s1;
  --sdram_0_s1_writedata mux, which is an e_mux
  sdram_0_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_nios2_clock_8_out_granted_sdram_0_s1)) = '1'), nios2_clock_8_out_writedata, nios2_clock_9_out_writedata);
  internal_nios2_clock_9_out_requests_sdram_0_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_9_out_read OR nios2_clock_9_out_write)))))));
  --nios2_clock_8/out granted sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_clock_8_out_granted_slave_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_clock_8_out_granted_slave_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_clock_8_out_saved_grant_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_0_s1_arbitration_holdoff_internal OR NOT internal_nios2_clock_8_out_requests_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_clock_8_out_granted_slave_sdram_0_s1))))));
    end if;

  end process;

  --nios2_clock_8_out_continuerequest continued request, which is an e_mux
  nios2_clock_8_out_continuerequest <= last_cycle_nios2_clock_8_out_granted_slave_sdram_0_s1 AND internal_nios2_clock_8_out_requests_sdram_0_s1;
  internal_nios2_clock_9_out_qualified_request_sdram_0_s1 <= internal_nios2_clock_9_out_requests_sdram_0_s1 AND NOT ((((nios2_clock_9_out_read AND (internal_nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register))) OR nios2_clock_8_out_arbiterlock));
  --rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1 : rdv_fifo_for_nios2_clock_9_out_to_sdram_0_s1_module
    port map(
      data_out => nios2_clock_9_out_rdv_fifo_output_from_sdram_0_s1,
      empty => open,
      fifo_contains_ones_n => nios2_clock_9_out_rdv_fifo_empty_sdram_0_s1,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_nios2_clock_9_out_granted_sdram_0_s1,
      read => sdram_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT sdram_0_s1_waits_for_read;

  internal_nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register <= NOT nios2_clock_9_out_rdv_fifo_empty_sdram_0_s1;
  --local readdatavalid nios2_clock_9_out_read_data_valid_sdram_0_s1, which is an e_mux
  nios2_clock_9_out_read_data_valid_sdram_0_s1 <= ((sdram_0_s1_readdatavalid_from_sa AND nios2_clock_9_out_rdv_fifo_output_from_sdram_0_s1)) AND NOT nios2_clock_9_out_rdv_fifo_empty_sdram_0_s1;
  --allow new arb cycle for sdram_0/s1, which is an e_assign
  sdram_0_s1_allow_new_arb_cycle <= NOT nios2_clock_8_out_arbiterlock AND NOT nios2_clock_9_out_arbiterlock;
  --nios2_clock_9/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  sdram_0_s1_master_qreq_vector(0) <= internal_nios2_clock_9_out_qualified_request_sdram_0_s1;
  --nios2_clock_9/out grant sdram_0/s1, which is an e_assign
  internal_nios2_clock_9_out_granted_sdram_0_s1 <= sdram_0_s1_grant_vector(0);
  --nios2_clock_9/out saved-grant sdram_0/s1, which is an e_assign
  nios2_clock_9_out_saved_grant_sdram_0_s1 <= sdram_0_s1_arb_winner(0) AND internal_nios2_clock_9_out_requests_sdram_0_s1;
  --nios2_clock_8/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  sdram_0_s1_master_qreq_vector(1) <= internal_nios2_clock_8_out_qualified_request_sdram_0_s1;
  --nios2_clock_8/out grant sdram_0/s1, which is an e_assign
  internal_nios2_clock_8_out_granted_sdram_0_s1 <= sdram_0_s1_grant_vector(1);
  --nios2_clock_8/out saved-grant sdram_0/s1, which is an e_assign
  nios2_clock_8_out_saved_grant_sdram_0_s1 <= sdram_0_s1_arb_winner(1) AND internal_nios2_clock_8_out_requests_sdram_0_s1;
  --sdram_0/s1 chosen-master double-vector, which is an e_assign
  sdram_0_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sdram_0_s1_master_qreq_vector & sdram_0_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sdram_0_s1_master_qreq_vector & NOT sdram_0_s1_master_qreq_vector))) + (std_logic_vector'("000") & (sdram_0_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  sdram_0_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((sdram_0_s1_allow_new_arb_cycle AND or_reduce(sdram_0_s1_grant_vector)))) = '1'), sdram_0_s1_grant_vector, sdram_0_s1_saved_chosen_master_vector);
  --saved sdram_0_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_0_s1_allow_new_arb_cycle) = '1' then 
        sdram_0_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sdram_0_s1_grant_vector)) = '1'), sdram_0_s1_grant_vector, sdram_0_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sdram_0_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sdram_0_s1_chosen_master_double_vector(1) OR sdram_0_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((sdram_0_s1_chosen_master_double_vector(0) OR sdram_0_s1_chosen_master_double_vector(2)))));
  --sdram_0/s1 chosen master rotated left, which is an e_assign
  sdram_0_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sdram_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(sdram_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --sdram_0/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sdram_0_s1_grant_vector)) = '1' then 
        sdram_0_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(sdram_0_s1_end_xfer) = '1'), sdram_0_s1_chosen_master_rot_left, sdram_0_s1_grant_vector);
      end if;
    end if;

  end process;

  --sdram_0_s1_reset_n assignment, which is an e_assign
  sdram_0_s1_reset_n <= reset_n;
  sdram_0_s1_chipselect <= internal_nios2_clock_8_out_granted_sdram_0_s1 OR internal_nios2_clock_9_out_granted_sdram_0_s1;
  --sdram_0_s1_firsttransfer first transaction, which is an e_assign
  sdram_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sdram_0_s1_begins_xfer) = '1'), sdram_0_s1_unreg_firsttransfer, sdram_0_s1_reg_firsttransfer);
  --sdram_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  sdram_0_s1_unreg_firsttransfer <= NOT ((sdram_0_s1_slavearbiterlockenable AND sdram_0_s1_any_continuerequest));
  --sdram_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_0_s1_begins_xfer) = '1' then 
        sdram_0_s1_reg_firsttransfer <= sdram_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sdram_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sdram_0_s1_beginbursttransfer_internal <= sdram_0_s1_begins_xfer;
  --sdram_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sdram_0_s1_arbitration_holdoff_internal <= sdram_0_s1_begins_xfer AND sdram_0_s1_firsttransfer;
  --~sdram_0_s1_read_n assignment, which is an e_mux
  sdram_0_s1_read_n <= NOT ((((internal_nios2_clock_8_out_granted_sdram_0_s1 AND nios2_clock_8_out_read)) OR ((internal_nios2_clock_9_out_granted_sdram_0_s1 AND nios2_clock_9_out_read))));
  --~sdram_0_s1_write_n assignment, which is an e_mux
  sdram_0_s1_write_n <= NOT ((((internal_nios2_clock_8_out_granted_sdram_0_s1 AND nios2_clock_8_out_write)) OR ((internal_nios2_clock_9_out_granted_sdram_0_s1 AND nios2_clock_9_out_write))));
  shifted_address_to_sdram_0_s1_from_nios2_clock_8_out <= nios2_clock_8_out_address_to_slave;
  --sdram_0_s1_address mux, which is an e_mux
  sdram_0_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_clock_8_out_granted_sdram_0_s1)) = '1'), (A_SRL(shifted_address_to_sdram_0_s1_from_nios2_clock_8_out,std_logic_vector'("00000000000000000000000000000001"))), (A_SRL(shifted_address_to_sdram_0_s1_from_nios2_clock_9_out,std_logic_vector'("00000000000000000000000000000001")))), 22);
  shifted_address_to_sdram_0_s1_from_nios2_clock_9_out <= nios2_clock_9_out_address_to_slave;
  --d1_sdram_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sdram_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sdram_0_s1_end_xfer <= sdram_0_s1_end_xfer;
    end if;

  end process;

  --sdram_0_s1_waits_for_read in a cycle, which is an e_mux
  sdram_0_s1_waits_for_read <= sdram_0_s1_in_a_read_cycle AND internal_sdram_0_s1_waitrequest_from_sa;
  --sdram_0_s1_in_a_read_cycle assignment, which is an e_assign
  sdram_0_s1_in_a_read_cycle <= ((internal_nios2_clock_8_out_granted_sdram_0_s1 AND nios2_clock_8_out_read)) OR ((internal_nios2_clock_9_out_granted_sdram_0_s1 AND nios2_clock_9_out_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sdram_0_s1_in_a_read_cycle;
  --sdram_0_s1_waits_for_write in a cycle, which is an e_mux
  sdram_0_s1_waits_for_write <= sdram_0_s1_in_a_write_cycle AND internal_sdram_0_s1_waitrequest_from_sa;
  --sdram_0_s1_in_a_write_cycle assignment, which is an e_assign
  sdram_0_s1_in_a_write_cycle <= ((internal_nios2_clock_8_out_granted_sdram_0_s1 AND nios2_clock_8_out_write)) OR ((internal_nios2_clock_9_out_granted_sdram_0_s1 AND nios2_clock_9_out_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sdram_0_s1_in_a_write_cycle;
  wait_for_sdram_0_s1_counter <= std_logic'('0');
  --~sdram_0_s1_byteenable_n byte enable port mux, which is an e_mux
  sdram_0_s1_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_nios2_clock_8_out_granted_sdram_0_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (nios2_clock_8_out_byteenable)), A_WE_StdLogicVector((std_logic'((internal_nios2_clock_9_out_granted_sdram_0_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (nios2_clock_9_out_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))), 2);
  --vhdl renameroo for output signals
  nios2_clock_8_out_granted_sdram_0_s1 <= internal_nios2_clock_8_out_granted_sdram_0_s1;
  --vhdl renameroo for output signals
  nios2_clock_8_out_qualified_request_sdram_0_s1 <= internal_nios2_clock_8_out_qualified_request_sdram_0_s1;
  --vhdl renameroo for output signals
  nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register <= internal_nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register;
  --vhdl renameroo for output signals
  nios2_clock_8_out_requests_sdram_0_s1 <= internal_nios2_clock_8_out_requests_sdram_0_s1;
  --vhdl renameroo for output signals
  nios2_clock_9_out_granted_sdram_0_s1 <= internal_nios2_clock_9_out_granted_sdram_0_s1;
  --vhdl renameroo for output signals
  nios2_clock_9_out_qualified_request_sdram_0_s1 <= internal_nios2_clock_9_out_qualified_request_sdram_0_s1;
  --vhdl renameroo for output signals
  nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register <= internal_nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register;
  --vhdl renameroo for output signals
  nios2_clock_9_out_requests_sdram_0_s1 <= internal_nios2_clock_9_out_requests_sdram_0_s1;
  --vhdl renameroo for output signals
  sdram_0_s1_waitrequest_from_sa <= internal_sdram_0_s1_waitrequest_from_sa;
--synthesis translate_off
    --sdram_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line99 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_clock_8_out_granted_sdram_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_clock_9_out_granted_sdram_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line99, now);
          write(write_line99, string'(": "));
          write(write_line99, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line99.all);
          deallocate (write_line99);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line100 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_clock_8_out_saved_grant_sdram_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_clock_9_out_saved_grant_sdram_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line100, now);
          write(write_line100, string'(": "));
          write(write_line100, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line100.all);
          deallocate (write_line100);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity switch_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_14_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_14_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_14_out_read : IN STD_LOGIC;
                 signal nios2_clock_14_out_write : IN STD_LOGIC;
                 signal nios2_clock_14_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal switch_pio_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- outputs:
                 signal d1_switch_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_14_out_granted_switch_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_14_out_qualified_request_switch_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_14_out_read_data_valid_switch_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_14_out_requests_switch_pio_s1 : OUT STD_LOGIC;
                 signal switch_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal switch_pio_s1_chipselect : OUT STD_LOGIC;
                 signal switch_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal switch_pio_s1_reset_n : OUT STD_LOGIC;
                 signal switch_pio_s1_write_n : OUT STD_LOGIC;
                 signal switch_pio_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
              );
end entity switch_pio_s1_arbitrator;


architecture europa of switch_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_switch_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_14_out_granted_switch_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_14_out_qualified_request_switch_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_14_out_requests_switch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_14_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_14_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_14_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_14_out_saved_grant_switch_pio_s1 :  STD_LOGIC;
                signal switch_pio_s1_allgrants :  STD_LOGIC;
                signal switch_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal switch_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal switch_pio_s1_any_continuerequest :  STD_LOGIC;
                signal switch_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal switch_pio_s1_arb_share_counter :  STD_LOGIC;
                signal switch_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal switch_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal switch_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal switch_pio_s1_begins_xfer :  STD_LOGIC;
                signal switch_pio_s1_end_xfer :  STD_LOGIC;
                signal switch_pio_s1_firsttransfer :  STD_LOGIC;
                signal switch_pio_s1_grant_vector :  STD_LOGIC;
                signal switch_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal switch_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal switch_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal switch_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal switch_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal switch_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal switch_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal switch_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal switch_pio_s1_waits_for_read :  STD_LOGIC;
                signal switch_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_switch_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT switch_pio_s1_end_xfer;
    end if;

  end process;

  switch_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_14_out_qualified_request_switch_pio_s1);
  --assign switch_pio_s1_readdata_from_sa = switch_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  switch_pio_s1_readdata_from_sa <= switch_pio_s1_readdata;
  internal_nios2_clock_14_out_requests_switch_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_14_out_read OR nios2_clock_14_out_write)))))));
  --switch_pio_s1_arb_share_counter set values, which is an e_mux
  switch_pio_s1_arb_share_set_values <= std_logic'('1');
  --switch_pio_s1_non_bursting_master_requests mux, which is an e_mux
  switch_pio_s1_non_bursting_master_requests <= internal_nios2_clock_14_out_requests_switch_pio_s1;
  --switch_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  switch_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --switch_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  switch_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(switch_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(switch_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(switch_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(switch_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --switch_pio_s1_allgrants all slave grants, which is an e_mux
  switch_pio_s1_allgrants <= switch_pio_s1_grant_vector;
  --switch_pio_s1_end_xfer assignment, which is an e_assign
  switch_pio_s1_end_xfer <= NOT ((switch_pio_s1_waits_for_read OR switch_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_switch_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_switch_pio_s1 <= switch_pio_s1_end_xfer AND (((NOT switch_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --switch_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  switch_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_switch_pio_s1 AND switch_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_switch_pio_s1 AND NOT switch_pio_s1_non_bursting_master_requests));
  --switch_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      switch_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(switch_pio_s1_arb_counter_enable) = '1' then 
        switch_pio_s1_arb_share_counter <= switch_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --switch_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      switch_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((switch_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_switch_pio_s1)) OR ((end_xfer_arb_share_counter_term_switch_pio_s1 AND NOT switch_pio_s1_non_bursting_master_requests)))) = '1' then 
        switch_pio_s1_slavearbiterlockenable <= switch_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_14/out switch_pio/s1 arbiterlock, which is an e_assign
  nios2_clock_14_out_arbiterlock <= switch_pio_s1_slavearbiterlockenable AND nios2_clock_14_out_continuerequest;
  --switch_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  switch_pio_s1_slavearbiterlockenable2 <= switch_pio_s1_arb_share_counter_next_value;
  --nios2_clock_14/out switch_pio/s1 arbiterlock2, which is an e_assign
  nios2_clock_14_out_arbiterlock2 <= switch_pio_s1_slavearbiterlockenable2 AND nios2_clock_14_out_continuerequest;
  --switch_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  switch_pio_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_14_out_continuerequest continued request, which is an e_assign
  nios2_clock_14_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_14_out_qualified_request_switch_pio_s1 <= internal_nios2_clock_14_out_requests_switch_pio_s1;
  --switch_pio_s1_writedata mux, which is an e_mux
  switch_pio_s1_writedata <= nios2_clock_14_out_writedata (3 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_clock_14_out_granted_switch_pio_s1 <= internal_nios2_clock_14_out_qualified_request_switch_pio_s1;
  --nios2_clock_14/out saved-grant switch_pio/s1, which is an e_assign
  nios2_clock_14_out_saved_grant_switch_pio_s1 <= internal_nios2_clock_14_out_requests_switch_pio_s1;
  --allow new arb cycle for switch_pio/s1, which is an e_assign
  switch_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  switch_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  switch_pio_s1_master_qreq_vector <= std_logic'('1');
  --switch_pio_s1_reset_n assignment, which is an e_assign
  switch_pio_s1_reset_n <= reset_n;
  switch_pio_s1_chipselect <= internal_nios2_clock_14_out_granted_switch_pio_s1;
  --switch_pio_s1_firsttransfer first transaction, which is an e_assign
  switch_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(switch_pio_s1_begins_xfer) = '1'), switch_pio_s1_unreg_firsttransfer, switch_pio_s1_reg_firsttransfer);
  --switch_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  switch_pio_s1_unreg_firsttransfer <= NOT ((switch_pio_s1_slavearbiterlockenable AND switch_pio_s1_any_continuerequest));
  --switch_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      switch_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(switch_pio_s1_begins_xfer) = '1' then 
        switch_pio_s1_reg_firsttransfer <= switch_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --switch_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  switch_pio_s1_beginbursttransfer_internal <= switch_pio_s1_begins_xfer;
  --~switch_pio_s1_write_n assignment, which is an e_mux
  switch_pio_s1_write_n <= NOT ((internal_nios2_clock_14_out_granted_switch_pio_s1 AND nios2_clock_14_out_write));
  --switch_pio_s1_address mux, which is an e_mux
  switch_pio_s1_address <= nios2_clock_14_out_nativeaddress;
  --d1_switch_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_switch_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_switch_pio_s1_end_xfer <= switch_pio_s1_end_xfer;
    end if;

  end process;

  --switch_pio_s1_waits_for_read in a cycle, which is an e_mux
  switch_pio_s1_waits_for_read <= switch_pio_s1_in_a_read_cycle AND switch_pio_s1_begins_xfer;
  --switch_pio_s1_in_a_read_cycle assignment, which is an e_assign
  switch_pio_s1_in_a_read_cycle <= internal_nios2_clock_14_out_granted_switch_pio_s1 AND nios2_clock_14_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= switch_pio_s1_in_a_read_cycle;
  --switch_pio_s1_waits_for_write in a cycle, which is an e_mux
  switch_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(switch_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --switch_pio_s1_in_a_write_cycle assignment, which is an e_assign
  switch_pio_s1_in_a_write_cycle <= internal_nios2_clock_14_out_granted_switch_pio_s1 AND nios2_clock_14_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= switch_pio_s1_in_a_write_cycle;
  wait_for_switch_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_14_out_granted_switch_pio_s1 <= internal_nios2_clock_14_out_granted_switch_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_14_out_qualified_request_switch_pio_s1 <= internal_nios2_clock_14_out_qualified_request_switch_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_14_out_requests_switch_pio_s1 <= internal_nios2_clock_14_out_requests_switch_pio_s1;
--synthesis translate_off
    --switch_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sys_clk_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_3_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_3_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_3_out_read : IN STD_LOGIC;
                 signal nios2_clock_3_out_write : IN STD_LOGIC;
                 signal nios2_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                 signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_3_out_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal nios2_clock_3_out_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal nios2_clock_3_out_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal nios2_clock_3_out_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sys_clk_timer_s1_arbitrator;


architecture europa of sys_clk_timer_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sys_clk_timer_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_3_out_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_nios2_clock_3_out_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_nios2_clock_3_out_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal nios2_clock_3_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_3_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_3_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_3_out_saved_grant_sys_clk_timer_s1 :  STD_LOGIC;
                signal sys_clk_timer_s1_allgrants :  STD_LOGIC;
                signal sys_clk_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sys_clk_timer_s1_any_continuerequest :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_counter :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_set_values :  STD_LOGIC;
                signal sys_clk_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sys_clk_timer_s1_begins_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_grant_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sys_clk_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sys_clk_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_read :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sys_clk_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  sys_clk_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_3_out_qualified_request_sys_clk_timer_s1);
  --assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_readdata_from_sa <= sys_clk_timer_s1_readdata;
  internal_nios2_clock_3_out_requests_sys_clk_timer_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_3_out_read OR nios2_clock_3_out_write)))))));
  --sys_clk_timer_s1_arb_share_counter set values, which is an e_mux
  sys_clk_timer_s1_arb_share_set_values <= std_logic'('1');
  --sys_clk_timer_s1_non_bursting_master_requests mux, which is an e_mux
  sys_clk_timer_s1_non_bursting_master_requests <= internal_nios2_clock_3_out_requests_sys_clk_timer_s1;
  --sys_clk_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sys_clk_timer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sys_clk_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  sys_clk_timer_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sys_clk_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sys_clk_timer_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sys_clk_timer_s1_allgrants all slave grants, which is an e_mux
  sys_clk_timer_s1_allgrants <= sys_clk_timer_s1_grant_vector;
  --sys_clk_timer_s1_end_xfer assignment, which is an e_assign
  sys_clk_timer_s1_end_xfer <= NOT ((sys_clk_timer_s1_waits_for_read OR sys_clk_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sys_clk_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sys_clk_timer_s1 <= sys_clk_timer_s1_end_xfer AND (((NOT sys_clk_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sys_clk_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sys_clk_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND sys_clk_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests));
  --sys_clk_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_arb_counter_enable) = '1' then 
        sys_clk_timer_s1_arb_share_counter <= sys_clk_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sys_clk_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sys_clk_timer_s1)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests)))) = '1' then 
        sys_clk_timer_s1_slavearbiterlockenable <= sys_clk_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_3/out sys_clk_timer/s1 arbiterlock, which is an e_assign
  nios2_clock_3_out_arbiterlock <= sys_clk_timer_s1_slavearbiterlockenable AND nios2_clock_3_out_continuerequest;
  --sys_clk_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sys_clk_timer_s1_slavearbiterlockenable2 <= sys_clk_timer_s1_arb_share_counter_next_value;
  --nios2_clock_3/out sys_clk_timer/s1 arbiterlock2, which is an e_assign
  nios2_clock_3_out_arbiterlock2 <= sys_clk_timer_s1_slavearbiterlockenable2 AND nios2_clock_3_out_continuerequest;
  --sys_clk_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sys_clk_timer_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_3_out_continuerequest continued request, which is an e_assign
  nios2_clock_3_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_3_out_qualified_request_sys_clk_timer_s1 <= internal_nios2_clock_3_out_requests_sys_clk_timer_s1;
  --sys_clk_timer_s1_writedata mux, which is an e_mux
  sys_clk_timer_s1_writedata <= nios2_clock_3_out_writedata;
  --master is always granted when requested
  internal_nios2_clock_3_out_granted_sys_clk_timer_s1 <= internal_nios2_clock_3_out_qualified_request_sys_clk_timer_s1;
  --nios2_clock_3/out saved-grant sys_clk_timer/s1, which is an e_assign
  nios2_clock_3_out_saved_grant_sys_clk_timer_s1 <= internal_nios2_clock_3_out_requests_sys_clk_timer_s1;
  --allow new arb cycle for sys_clk_timer/s1, which is an e_assign
  sys_clk_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sys_clk_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sys_clk_timer_s1_master_qreq_vector <= std_logic'('1');
  --sys_clk_timer_s1_reset_n assignment, which is an e_assign
  sys_clk_timer_s1_reset_n <= reset_n;
  sys_clk_timer_s1_chipselect <= internal_nios2_clock_3_out_granted_sys_clk_timer_s1;
  --sys_clk_timer_s1_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sys_clk_timer_s1_begins_xfer) = '1'), sys_clk_timer_s1_unreg_firsttransfer, sys_clk_timer_s1_reg_firsttransfer);
  --sys_clk_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_unreg_firsttransfer <= NOT ((sys_clk_timer_s1_slavearbiterlockenable AND sys_clk_timer_s1_any_continuerequest));
  --sys_clk_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_begins_xfer) = '1' then 
        sys_clk_timer_s1_reg_firsttransfer <= sys_clk_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sys_clk_timer_s1_beginbursttransfer_internal <= sys_clk_timer_s1_begins_xfer;
  --~sys_clk_timer_s1_write_n assignment, which is an e_mux
  sys_clk_timer_s1_write_n <= NOT ((internal_nios2_clock_3_out_granted_sys_clk_timer_s1 AND nios2_clock_3_out_write));
  --sys_clk_timer_s1_address mux, which is an e_mux
  sys_clk_timer_s1_address <= nios2_clock_3_out_nativeaddress;
  --d1_sys_clk_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sys_clk_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sys_clk_timer_s1_end_xfer <= sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  --sys_clk_timer_s1_waits_for_read in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_read <= sys_clk_timer_s1_in_a_read_cycle AND sys_clk_timer_s1_begins_xfer;
  --sys_clk_timer_s1_in_a_read_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_read_cycle <= internal_nios2_clock_3_out_granted_sys_clk_timer_s1 AND nios2_clock_3_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sys_clk_timer_s1_in_a_read_cycle;
  --sys_clk_timer_s1_waits_for_write in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sys_clk_timer_s1_in_a_write_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_write_cycle <= internal_nios2_clock_3_out_granted_sys_clk_timer_s1 AND nios2_clock_3_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sys_clk_timer_s1_in_a_write_cycle;
  wait_for_sys_clk_timer_s1_counter <= std_logic'('0');
  --assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_irq_from_sa <= sys_clk_timer_s1_irq;
  --vhdl renameroo for output signals
  nios2_clock_3_out_granted_sys_clk_timer_s1 <= internal_nios2_clock_3_out_granted_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  nios2_clock_3_out_qualified_request_sys_clk_timer_s1 <= internal_nios2_clock_3_out_qualified_request_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  nios2_clock_3_out_requests_sys_clk_timer_s1 <= internal_nios2_clock_3_out_requests_sys_clk_timer_s1;
--synthesis translate_off
    --sys_clk_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sysid_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_4_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_clock_4_out_nativeaddress : IN STD_LOGIC;
                 signal nios2_clock_4_out_read : IN STD_LOGIC;
                 signal nios2_clock_4_out_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_4_out_granted_sysid_control_slave : OUT STD_LOGIC;
                 signal nios2_clock_4_out_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                 signal nios2_clock_4_out_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                 signal nios2_clock_4_out_requests_sysid_control_slave : OUT STD_LOGIC;
                 signal sysid_control_slave_address : OUT STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sysid_control_slave_reset_n : OUT STD_LOGIC
              );
end entity sysid_control_slave_arbitrator;


architecture europa of sysid_control_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sysid_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_4_out_granted_sysid_control_slave :  STD_LOGIC;
                signal internal_nios2_clock_4_out_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal internal_nios2_clock_4_out_requests_sysid_control_slave :  STD_LOGIC;
                signal nios2_clock_4_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_4_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_4_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_4_out_saved_grant_sysid_control_slave :  STD_LOGIC;
                signal sysid_control_slave_allgrants :  STD_LOGIC;
                signal sysid_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal sysid_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sysid_control_slave_any_continuerequest :  STD_LOGIC;
                signal sysid_control_slave_arb_counter_enable :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal sysid_control_slave_arb_share_set_values :  STD_LOGIC;
                signal sysid_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal sysid_control_slave_begins_xfer :  STD_LOGIC;
                signal sysid_control_slave_end_xfer :  STD_LOGIC;
                signal sysid_control_slave_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_grant_vector :  STD_LOGIC;
                signal sysid_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal sysid_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal sysid_control_slave_master_qreq_vector :  STD_LOGIC;
                signal sysid_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal sysid_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal sysid_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_waits_for_read :  STD_LOGIC;
                signal sysid_control_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_sysid_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sysid_control_slave_end_xfer;
    end if;

  end process;

  sysid_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_4_out_qualified_request_sysid_control_slave);
  --assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysid_control_slave_readdata_from_sa <= sysid_control_slave_readdata;
  internal_nios2_clock_4_out_requests_sysid_control_slave <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_4_out_read OR nios2_clock_4_out_write))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_clock_4_out_read)))));
  --sysid_control_slave_arb_share_counter set values, which is an e_mux
  sysid_control_slave_arb_share_set_values <= std_logic'('1');
  --sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  sysid_control_slave_non_bursting_master_requests <= internal_nios2_clock_4_out_requests_sysid_control_slave;
  --sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  sysid_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  sysid_control_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sysid_control_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sysid_control_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sysid_control_slave_allgrants all slave grants, which is an e_mux
  sysid_control_slave_allgrants <= sysid_control_slave_grant_vector;
  --sysid_control_slave_end_xfer assignment, which is an e_assign
  sysid_control_slave_end_xfer <= NOT ((sysid_control_slave_waits_for_read OR sysid_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sysid_control_slave <= sysid_control_slave_end_xfer AND (((NOT sysid_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  sysid_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sysid_control_slave AND sysid_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests));
  --sysid_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_arb_counter_enable) = '1' then 
        sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sysid_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_sysid_control_slave)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests)))) = '1' then 
        sysid_control_slave_slavearbiterlockenable <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_4/out sysid/control_slave arbiterlock, which is an e_assign
  nios2_clock_4_out_arbiterlock <= sysid_control_slave_slavearbiterlockenable AND nios2_clock_4_out_continuerequest;
  --sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sysid_control_slave_slavearbiterlockenable2 <= sysid_control_slave_arb_share_counter_next_value;
  --nios2_clock_4/out sysid/control_slave arbiterlock2, which is an e_assign
  nios2_clock_4_out_arbiterlock2 <= sysid_control_slave_slavearbiterlockenable2 AND nios2_clock_4_out_continuerequest;
  --sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  sysid_control_slave_any_continuerequest <= std_logic'('1');
  --nios2_clock_4_out_continuerequest continued request, which is an e_assign
  nios2_clock_4_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_4_out_qualified_request_sysid_control_slave <= internal_nios2_clock_4_out_requests_sysid_control_slave;
  --master is always granted when requested
  internal_nios2_clock_4_out_granted_sysid_control_slave <= internal_nios2_clock_4_out_qualified_request_sysid_control_slave;
  --nios2_clock_4/out saved-grant sysid/control_slave, which is an e_assign
  nios2_clock_4_out_saved_grant_sysid_control_slave <= internal_nios2_clock_4_out_requests_sysid_control_slave;
  --allow new arb cycle for sysid/control_slave, which is an e_assign
  sysid_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sysid_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sysid_control_slave_master_qreq_vector <= std_logic'('1');
  --sysid_control_slave_reset_n assignment, which is an e_assign
  sysid_control_slave_reset_n <= reset_n;
  --sysid_control_slave_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(sysid_control_slave_begins_xfer) = '1'), sysid_control_slave_unreg_firsttransfer, sysid_control_slave_reg_firsttransfer);
  --sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_unreg_firsttransfer <= NOT ((sysid_control_slave_slavearbiterlockenable AND sysid_control_slave_any_continuerequest));
  --sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_begins_xfer) = '1' then 
        sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sysid_control_slave_beginbursttransfer_internal <= sysid_control_slave_begins_xfer;
  --sysid_control_slave_address mux, which is an e_mux
  sysid_control_slave_address <= nios2_clock_4_out_nativeaddress;
  --d1_sysid_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sysid_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end if;

  end process;

  --sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  sysid_control_slave_waits_for_read <= sysid_control_slave_in_a_read_cycle AND sysid_control_slave_begins_xfer;
  --sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_read_cycle <= internal_nios2_clock_4_out_granted_sysid_control_slave AND nios2_clock_4_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sysid_control_slave_in_a_read_cycle;
  --sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  sysid_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_write_cycle <= internal_nios2_clock_4_out_granted_sysid_control_slave AND nios2_clock_4_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sysid_control_slave_in_a_write_cycle;
  wait_for_sysid_control_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_4_out_granted_sysid_control_slave <= internal_nios2_clock_4_out_granted_sysid_control_slave;
  --vhdl renameroo for output signals
  nios2_clock_4_out_qualified_request_sysid_control_slave <= internal_nios2_clock_4_out_qualified_request_sysid_control_slave;
  --vhdl renameroo for output signals
  nios2_clock_4_out_requests_sysid_control_slave <= internal_nios2_clock_4_out_requests_sysid_control_slave;
--synthesis translate_off
    --sysid/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity usb_code_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_clock_16_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_clock_16_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_clock_16_out_read : IN STD_LOGIC;
                 signal nios2_clock_16_out_write : IN STD_LOGIC;
                 signal nios2_clock_16_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal usb_code_pio_s1_readdata : IN STD_LOGIC_VECTOR (20 DOWNTO 0);

              -- outputs:
                 signal d1_usb_code_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_clock_16_out_granted_usb_code_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_16_out_qualified_request_usb_code_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_16_out_read_data_valid_usb_code_pio_s1 : OUT STD_LOGIC;
                 signal nios2_clock_16_out_requests_usb_code_pio_s1 : OUT STD_LOGIC;
                 signal usb_code_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal usb_code_pio_s1_chipselect : OUT STD_LOGIC;
                 signal usb_code_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal usb_code_pio_s1_reset_n : OUT STD_LOGIC;
                 signal usb_code_pio_s1_write_n : OUT STD_LOGIC;
                 signal usb_code_pio_s1_writedata : OUT STD_LOGIC_VECTOR (20 DOWNTO 0)
              );
end entity usb_code_pio_s1_arbitrator;


architecture europa of usb_code_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_usb_code_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_clock_16_out_granted_usb_code_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_16_out_qualified_request_usb_code_pio_s1 :  STD_LOGIC;
                signal internal_nios2_clock_16_out_requests_usb_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_16_out_arbiterlock :  STD_LOGIC;
                signal nios2_clock_16_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_clock_16_out_continuerequest :  STD_LOGIC;
                signal nios2_clock_16_out_saved_grant_usb_code_pio_s1 :  STD_LOGIC;
                signal usb_code_pio_s1_allgrants :  STD_LOGIC;
                signal usb_code_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal usb_code_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal usb_code_pio_s1_any_continuerequest :  STD_LOGIC;
                signal usb_code_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal usb_code_pio_s1_arb_share_counter :  STD_LOGIC;
                signal usb_code_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal usb_code_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal usb_code_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal usb_code_pio_s1_begins_xfer :  STD_LOGIC;
                signal usb_code_pio_s1_end_xfer :  STD_LOGIC;
                signal usb_code_pio_s1_firsttransfer :  STD_LOGIC;
                signal usb_code_pio_s1_grant_vector :  STD_LOGIC;
                signal usb_code_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal usb_code_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal usb_code_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal usb_code_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal usb_code_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal usb_code_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal usb_code_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal usb_code_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal usb_code_pio_s1_waits_for_read :  STD_LOGIC;
                signal usb_code_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_usb_code_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT usb_code_pio_s1_end_xfer;
    end if;

  end process;

  usb_code_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_clock_16_out_qualified_request_usb_code_pio_s1);
  --assign usb_code_pio_s1_readdata_from_sa = usb_code_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  usb_code_pio_s1_readdata_from_sa <= usb_code_pio_s1_readdata;
  internal_nios2_clock_16_out_requests_usb_code_pio_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_clock_16_out_read OR nios2_clock_16_out_write)))))));
  --usb_code_pio_s1_arb_share_counter set values, which is an e_mux
  usb_code_pio_s1_arb_share_set_values <= std_logic'('1');
  --usb_code_pio_s1_non_bursting_master_requests mux, which is an e_mux
  usb_code_pio_s1_non_bursting_master_requests <= internal_nios2_clock_16_out_requests_usb_code_pio_s1;
  --usb_code_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  usb_code_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --usb_code_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  usb_code_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(usb_code_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(usb_code_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(usb_code_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(usb_code_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --usb_code_pio_s1_allgrants all slave grants, which is an e_mux
  usb_code_pio_s1_allgrants <= usb_code_pio_s1_grant_vector;
  --usb_code_pio_s1_end_xfer assignment, which is an e_assign
  usb_code_pio_s1_end_xfer <= NOT ((usb_code_pio_s1_waits_for_read OR usb_code_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_usb_code_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_usb_code_pio_s1 <= usb_code_pio_s1_end_xfer AND (((NOT usb_code_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --usb_code_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  usb_code_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_usb_code_pio_s1 AND usb_code_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_usb_code_pio_s1 AND NOT usb_code_pio_s1_non_bursting_master_requests));
  --usb_code_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      usb_code_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(usb_code_pio_s1_arb_counter_enable) = '1' then 
        usb_code_pio_s1_arb_share_counter <= usb_code_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --usb_code_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      usb_code_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((usb_code_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_usb_code_pio_s1)) OR ((end_xfer_arb_share_counter_term_usb_code_pio_s1 AND NOT usb_code_pio_s1_non_bursting_master_requests)))) = '1' then 
        usb_code_pio_s1_slavearbiterlockenable <= usb_code_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_clock_16/out usb_code_pio/s1 arbiterlock, which is an e_assign
  nios2_clock_16_out_arbiterlock <= usb_code_pio_s1_slavearbiterlockenable AND nios2_clock_16_out_continuerequest;
  --usb_code_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  usb_code_pio_s1_slavearbiterlockenable2 <= usb_code_pio_s1_arb_share_counter_next_value;
  --nios2_clock_16/out usb_code_pio/s1 arbiterlock2, which is an e_assign
  nios2_clock_16_out_arbiterlock2 <= usb_code_pio_s1_slavearbiterlockenable2 AND nios2_clock_16_out_continuerequest;
  --usb_code_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  usb_code_pio_s1_any_continuerequest <= std_logic'('1');
  --nios2_clock_16_out_continuerequest continued request, which is an e_assign
  nios2_clock_16_out_continuerequest <= std_logic'('1');
  internal_nios2_clock_16_out_qualified_request_usb_code_pio_s1 <= internal_nios2_clock_16_out_requests_usb_code_pio_s1;
  --usb_code_pio_s1_writedata mux, which is an e_mux
  usb_code_pio_s1_writedata <= nios2_clock_16_out_writedata (20 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_clock_16_out_granted_usb_code_pio_s1 <= internal_nios2_clock_16_out_qualified_request_usb_code_pio_s1;
  --nios2_clock_16/out saved-grant usb_code_pio/s1, which is an e_assign
  nios2_clock_16_out_saved_grant_usb_code_pio_s1 <= internal_nios2_clock_16_out_requests_usb_code_pio_s1;
  --allow new arb cycle for usb_code_pio/s1, which is an e_assign
  usb_code_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  usb_code_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  usb_code_pio_s1_master_qreq_vector <= std_logic'('1');
  --usb_code_pio_s1_reset_n assignment, which is an e_assign
  usb_code_pio_s1_reset_n <= reset_n;
  usb_code_pio_s1_chipselect <= internal_nios2_clock_16_out_granted_usb_code_pio_s1;
  --usb_code_pio_s1_firsttransfer first transaction, which is an e_assign
  usb_code_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(usb_code_pio_s1_begins_xfer) = '1'), usb_code_pio_s1_unreg_firsttransfer, usb_code_pio_s1_reg_firsttransfer);
  --usb_code_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  usb_code_pio_s1_unreg_firsttransfer <= NOT ((usb_code_pio_s1_slavearbiterlockenable AND usb_code_pio_s1_any_continuerequest));
  --usb_code_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      usb_code_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(usb_code_pio_s1_begins_xfer) = '1' then 
        usb_code_pio_s1_reg_firsttransfer <= usb_code_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --usb_code_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  usb_code_pio_s1_beginbursttransfer_internal <= usb_code_pio_s1_begins_xfer;
  --~usb_code_pio_s1_write_n assignment, which is an e_mux
  usb_code_pio_s1_write_n <= NOT ((internal_nios2_clock_16_out_granted_usb_code_pio_s1 AND nios2_clock_16_out_write));
  --usb_code_pio_s1_address mux, which is an e_mux
  usb_code_pio_s1_address <= nios2_clock_16_out_nativeaddress;
  --d1_usb_code_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_usb_code_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_usb_code_pio_s1_end_xfer <= usb_code_pio_s1_end_xfer;
    end if;

  end process;

  --usb_code_pio_s1_waits_for_read in a cycle, which is an e_mux
  usb_code_pio_s1_waits_for_read <= usb_code_pio_s1_in_a_read_cycle AND usb_code_pio_s1_begins_xfer;
  --usb_code_pio_s1_in_a_read_cycle assignment, which is an e_assign
  usb_code_pio_s1_in_a_read_cycle <= internal_nios2_clock_16_out_granted_usb_code_pio_s1 AND nios2_clock_16_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= usb_code_pio_s1_in_a_read_cycle;
  --usb_code_pio_s1_waits_for_write in a cycle, which is an e_mux
  usb_code_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(usb_code_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --usb_code_pio_s1_in_a_write_cycle assignment, which is an e_assign
  usb_code_pio_s1_in_a_write_cycle <= internal_nios2_clock_16_out_granted_usb_code_pio_s1 AND nios2_clock_16_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= usb_code_pio_s1_in_a_write_cycle;
  wait_for_usb_code_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_clock_16_out_granted_usb_code_pio_s1 <= internal_nios2_clock_16_out_granted_usb_code_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_16_out_qualified_request_usb_code_pio_s1 <= internal_nios2_clock_16_out_qualified_request_usb_code_pio_s1;
  --vhdl renameroo for output signals
  nios2_clock_16_out_requests_usb_code_pio_s1 <= internal_nios2_clock_16_out_requests_usb_code_pio_s1;
--synthesis translate_off
    --usb_code_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_reset_clk_0_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios2_reset_clk_0_domain_synch_module;


architecture europa of nios2_reset_clk_0_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_reset_altpll_0_c0_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios2_reset_altpll_0_c0_domain_synch_module;


architecture europa of nios2_reset_altpll_0_c0_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_reset_processor_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios2_reset_processor_clk_domain_synch_module;


architecture europa of nios2_reset_processor_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_reset_altpll_0_c1_out_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios2_reset_altpll_0_c1_out_domain_synch_module;


architecture europa of nios2_reset_altpll_0_c1_out_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2 is 
        port (
              -- 1) global signals:
                 signal altpll_0_c0 : OUT STD_LOGIC;
                 signal altpll_0_c1_out : OUT STD_LOGIC;
                 signal clk_0 : IN STD_LOGIC;
                 signal processor_clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- the_altpll_0
                 signal locked_from_the_altpll_0 : OUT STD_LOGIC;
                 signal phasedone_from_the_altpll_0 : OUT STD_LOGIC;

              -- the_cal_dac_code_pio
                 signal out_port_from_the_cal_dac_code_pio : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);

              -- the_comparator_pio
                 signal in_port_to_the_comparator_pio : IN STD_LOGIC;

              -- the_gen_code_strobe
                 signal out_port_from_the_gen_code_strobe : OUT STD_LOGIC;

              -- the_gen_code_value_pio_0
                 signal out_port_from_the_gen_code_value_pio_0 : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);

              -- the_gen_code_value_pio_1
                 signal out_port_from_the_gen_code_value_pio_1 : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);

              -- the_latch_pio
                 signal out_port_from_the_latch_pio : OUT STD_LOGIC;

              -- the_led_pio
                 signal out_port_from_the_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_mode_select
                 signal in_port_to_the_mode_select : IN STD_LOGIC_VECTOR (1 DOWNTO 0);

              -- the_sample_and_hold_pio
                 signal out_port_from_the_sample_and_hold_pio : OUT STD_LOGIC;

              -- the_sdram_0
                 signal zs_addr_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal zs_ba_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_cas_n_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_cke_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_cs_n_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_dq_to_and_from_the_sdram_0 : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal zs_dqm_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_ras_n_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_we_n_from_the_sdram_0 : OUT STD_LOGIC;

              -- the_switch_pio
                 signal out_port_from_the_switch_pio : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_usb_code_pio
                 signal out_port_from_the_usb_code_pio : OUT STD_LOGIC_VECTOR (20 DOWNTO 0)
              );
end entity nios2;


architecture europa of nios2 is
component altpll_0_pll_slave_arbitrator is 
           port (
                 -- inputs:
                    signal altpll_0_pll_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_5_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_5_out_read : IN STD_LOGIC;
                    signal nios2_clock_5_out_write : IN STD_LOGIC;
                    signal nios2_clock_5_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal altpll_0_pll_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal altpll_0_pll_slave_read : OUT STD_LOGIC;
                    signal altpll_0_pll_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal altpll_0_pll_slave_reset : OUT STD_LOGIC;
                    signal altpll_0_pll_slave_write : OUT STD_LOGIC;
                    signal altpll_0_pll_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_altpll_0_pll_slave_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_5_out_granted_altpll_0_pll_slave : OUT STD_LOGIC;
                    signal nios2_clock_5_out_qualified_request_altpll_0_pll_slave : OUT STD_LOGIC;
                    signal nios2_clock_5_out_read_data_valid_altpll_0_pll_slave : OUT STD_LOGIC;
                    signal nios2_clock_5_out_requests_altpll_0_pll_slave : OUT STD_LOGIC
                 );
end component altpll_0_pll_slave_arbitrator;

component altpll_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal c0 : OUT STD_LOGIC;
                    signal c1 : OUT STD_LOGIC;
                    signal locked : OUT STD_LOGIC;
                    signal phasedone : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component altpll_0;

component cal_dac_code_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal cal_dac_code_pio_s1_readdata : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_15_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_15_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_15_out_read : IN STD_LOGIC;
                    signal nios2_clock_15_out_write : IN STD_LOGIC;
                    signal nios2_clock_15_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cal_dac_code_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cal_dac_code_pio_s1_chipselect : OUT STD_LOGIC;
                    signal cal_dac_code_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal cal_dac_code_pio_s1_reset_n : OUT STD_LOGIC;
                    signal cal_dac_code_pio_s1_write_n : OUT STD_LOGIC;
                    signal cal_dac_code_pio_s1_writedata : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal d1_cal_dac_code_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_15_out_granted_cal_dac_code_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_15_out_requests_cal_dac_code_pio_s1 : OUT STD_LOGIC
                 );
end component cal_dac_code_pio_s1_arbitrator;

component cal_dac_code_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (13 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (13 DOWNTO 0)
                 );
end component cal_dac_code_pio;

component comparator_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal comparator_pio_s1_readdata : IN STD_LOGIC;
                    signal nios2_clock_11_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_11_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_11_out_read : IN STD_LOGIC;
                    signal nios2_clock_11_out_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal comparator_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal comparator_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal comparator_pio_s1_reset_n : OUT STD_LOGIC;
                    signal d1_comparator_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_11_out_granted_comparator_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_11_out_qualified_request_comparator_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_11_out_read_data_valid_comparator_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_11_out_requests_comparator_pio_s1 : OUT STD_LOGIC
                 );
end component comparator_pio_s1_arbitrator;

component comparator_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC
                 );
end component comparator_pio;

component cpu_0_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal cpu_0_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_reset_n : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_write : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_0_jtag_debug_module_end_xfer : OUT STD_LOGIC
                 );
end component cpu_0_jtag_debug_module_arbitrator;

component cpu_0_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_byteenable_nios2_clock_9_in : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_10_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_11_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_12_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_13_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_14_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_15_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_16_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_17_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_18_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_2_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_3_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_4_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_5_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_6_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_7_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_nios2_clock_9_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_10_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_11_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_12_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_13_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_14_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_15_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_16_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_17_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_18_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_2_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_3_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_4_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_5_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_6_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_7_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_9_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_10_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_11_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_12_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_13_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_14_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_15_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_16_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_17_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_18_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_2_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_3_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_4_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_5_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_6_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_7_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_9_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_10_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_11_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_12_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_13_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_14_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_15_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_16_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_17_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_18_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_2_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_3_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_4_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_5_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_6_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_7_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_9_in : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_10_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_11_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_12_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_13_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_14_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_15_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_16_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_17_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_18_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_1_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_2_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_3_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_4_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_5_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_6_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_7_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_9_in_end_xfer : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal nios2_clock_10_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_10_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_11_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_11_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_12_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_12_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_13_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_13_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_14_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_14_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_15_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_15_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_16_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_16_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_17_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_17_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_18_in_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_18_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_2_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_2_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_3_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_3_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_4_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_4_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_5_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_5_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_6_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_6_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_7_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_7_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_9_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_9_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal processor_clk : IN STD_LOGIC;
                    signal processor_clk_reset_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_0_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_0_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : OUT STD_LOGIC;
                    signal cpu_0_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_data_master_readdatavalid : OUT STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_0_data_master_arbitrator;

component cpu_0_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_instruction_master_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_granted_nios2_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_instruction_master_granted_nios2_clock_8_in : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_nios2_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_nios2_clock_8_in : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_nios2_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_nios2_clock_8_in : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_nios2_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_nios2_clock_8_in : IN STD_LOGIC;
                    signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_0_in_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_clock_8_in_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_8_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_8_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_0_instruction_master_latency_counter : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_0_instruction_master_arbitrator;

component cpu_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdatavalid : IN STD_LOGIC;
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component cpu_0;

component gen_code_strobe_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal gen_code_strobe_s1_readdata : IN STD_LOGIC;
                    signal nios2_clock_13_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_13_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_13_out_read : IN STD_LOGIC;
                    signal nios2_clock_13_out_write : IN STD_LOGIC;
                    signal nios2_clock_13_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_gen_code_strobe_s1_end_xfer : OUT STD_LOGIC;
                    signal gen_code_strobe_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gen_code_strobe_s1_chipselect : OUT STD_LOGIC;
                    signal gen_code_strobe_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal gen_code_strobe_s1_reset_n : OUT STD_LOGIC;
                    signal gen_code_strobe_s1_write_n : OUT STD_LOGIC;
                    signal gen_code_strobe_s1_writedata : OUT STD_LOGIC;
                    signal nios2_clock_13_out_granted_gen_code_strobe_s1 : OUT STD_LOGIC;
                    signal nios2_clock_13_out_qualified_request_gen_code_strobe_s1 : OUT STD_LOGIC;
                    signal nios2_clock_13_out_read_data_valid_gen_code_strobe_s1 : OUT STD_LOGIC;
                    signal nios2_clock_13_out_requests_gen_code_strobe_s1 : OUT STD_LOGIC
                 );
end component gen_code_strobe_s1_arbitrator;

component gen_code_strobe is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component gen_code_strobe;

component gen_code_value_pio_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal gen_code_value_pio_0_s1_readdata : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal nios2_clock_6_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_6_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_6_out_read : IN STD_LOGIC;
                    signal nios2_clock_6_out_write : IN STD_LOGIC;
                    signal nios2_clock_6_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_gen_code_value_pio_0_s1_end_xfer : OUT STD_LOGIC;
                    signal gen_code_value_pio_0_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gen_code_value_pio_0_s1_chipselect : OUT STD_LOGIC;
                    signal gen_code_value_pio_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal gen_code_value_pio_0_s1_reset_n : OUT STD_LOGIC;
                    signal gen_code_value_pio_0_s1_write_n : OUT STD_LOGIC;
                    signal gen_code_value_pio_0_s1_writedata : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal nios2_clock_6_out_granted_gen_code_value_pio_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_6_out_requests_gen_code_value_pio_0_s1 : OUT STD_LOGIC
                 );
end component gen_code_value_pio_0_s1_arbitrator;

component gen_code_value_pio_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (23 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (23 DOWNTO 0)
                 );
end component gen_code_value_pio_0;

component gen_code_value_pio_1_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal gen_code_value_pio_1_s1_readdata : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal nios2_clock_7_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_7_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_7_out_read : IN STD_LOGIC;
                    signal nios2_clock_7_out_write : IN STD_LOGIC;
                    signal nios2_clock_7_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_gen_code_value_pio_1_s1_end_xfer : OUT STD_LOGIC;
                    signal gen_code_value_pio_1_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gen_code_value_pio_1_s1_chipselect : OUT STD_LOGIC;
                    signal gen_code_value_pio_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal gen_code_value_pio_1_s1_reset_n : OUT STD_LOGIC;
                    signal gen_code_value_pio_1_s1_write_n : OUT STD_LOGIC;
                    signal gen_code_value_pio_1_s1_writedata : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal nios2_clock_7_out_granted_gen_code_value_pio_1_s1 : OUT STD_LOGIC;
                    signal nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 : OUT STD_LOGIC;
                    signal nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1 : OUT STD_LOGIC;
                    signal nios2_clock_7_out_requests_gen_code_value_pio_1_s1 : OUT STD_LOGIC
                 );
end component gen_code_value_pio_1_s1_arbitrator;

component gen_code_value_pio_1 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (23 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (23 DOWNTO 0)
                 );
end component gen_code_value_pio_1;

component jtag_uart_0_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_0_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal nios2_clock_2_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_2_out_nativeaddress : IN STD_LOGIC;
                    signal nios2_clock_2_out_read : IN STD_LOGIC;
                    signal nios2_clock_2_out_write : IN STD_LOGIC;
                    signal nios2_clock_2_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                    signal nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                    signal nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                    signal nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC
                 );
end component jtag_uart_0_avalon_jtag_slave_arbitrator;

component jtag_uart_0 is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart_0;

component latch_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal latch_pio_s1_readdata : IN STD_LOGIC;
                    signal nios2_clock_18_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_18_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_18_out_read : IN STD_LOGIC;
                    signal nios2_clock_18_out_write : IN STD_LOGIC;
                    signal nios2_clock_18_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_latch_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal latch_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal latch_pio_s1_chipselect : OUT STD_LOGIC;
                    signal latch_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal latch_pio_s1_reset_n : OUT STD_LOGIC;
                    signal latch_pio_s1_write_n : OUT STD_LOGIC;
                    signal latch_pio_s1_writedata : OUT STD_LOGIC;
                    signal nios2_clock_18_out_granted_latch_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_18_out_qualified_request_latch_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_18_out_read_data_valid_latch_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_18_out_requests_latch_pio_s1 : OUT STD_LOGIC
                 );
end component latch_pio_s1_arbitrator;

component latch_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component latch_pio;

component led_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_12_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_12_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_12_out_read : IN STD_LOGIC;
                    signal nios2_clock_12_out_write : IN STD_LOGIC;
                    signal nios2_clock_12_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal led_pio_s1_chipselect : OUT STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal led_pio_s1_reset_n : OUT STD_LOGIC;
                    signal led_pio_s1_write_n : OUT STD_LOGIC;
                    signal led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_12_out_granted_led_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_12_out_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_12_out_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_12_out_requests_led_pio_s1 : OUT STD_LOGIC
                 );
end component led_pio_s1_arbitrator;

component led_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component led_pio;

component mode_select_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal mode_select_s1_readdata : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_out_read : IN STD_LOGIC;
                    signal nios2_clock_10_out_write : IN STD_LOGIC;
                    signal nios2_clock_10_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_mode_select_s1_end_xfer : OUT STD_LOGIC;
                    signal mode_select_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mode_select_s1_chipselect : OUT STD_LOGIC;
                    signal mode_select_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mode_select_s1_reset_n : OUT STD_LOGIC;
                    signal mode_select_s1_write_n : OUT STD_LOGIC;
                    signal mode_select_s1_writedata : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_out_granted_mode_select_s1 : OUT STD_LOGIC;
                    signal nios2_clock_10_out_qualified_request_mode_select_s1 : OUT STD_LOGIC;
                    signal nios2_clock_10_out_read_data_valid_mode_select_s1 : OUT STD_LOGIC;
                    signal nios2_clock_10_out_requests_mode_select_s1 : OUT STD_LOGIC
                 );
end component mode_select_s1_arbitrator;

component mode_select is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (1 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
                 );
end component mode_select;

component nios2_clock_0_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal nios2_clock_0_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_0_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_instruction_master_granted_nios2_clock_0_in : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_nios2_clock_0_in : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_nios2_clock_0_in : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_nios2_clock_0_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_0_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_0_in_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_clock_0_in_read : OUT STD_LOGIC;
                    signal nios2_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_0_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_0_in_write : OUT STD_LOGIC
                 );
end component nios2_clock_0_in_arbitrator;

component nios2_clock_0_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_onchip_mem_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_0_out_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_0_out_granted_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_0_out_qualified_request_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_0_out_read : IN STD_LOGIC;
                    signal nios2_clock_0_out_read_data_valid_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_0_out_requests_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_0_out_write : IN STD_LOGIC;
                    signal nios2_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal onchip_mem_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_0_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_0_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_0_out_arbitrator;

component nios2_clock_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_0;

component nios2_clock_1_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_1_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_1_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_1_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_1_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_1_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_1_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_1_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_1_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_1_in_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_1_in_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_clock_1_in_read : OUT STD_LOGIC;
                    signal nios2_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_1_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_1_in_write : OUT STD_LOGIC;
                    signal nios2_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_clock_1_in_arbitrator;

component nios2_clock_1_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_onchip_mem_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_1_out_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_1_out_granted_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_1_out_qualified_request_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_1_out_read : IN STD_LOGIC;
                    signal nios2_clock_1_out_read_data_valid_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_1_out_requests_onchip_mem_s1 : IN STD_LOGIC;
                    signal nios2_clock_1_out_write : IN STD_LOGIC;
                    signal nios2_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal onchip_mem_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_1_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_1_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_1_out_arbitrator;

component nios2_clock_1 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_1;

component nios2_clock_10_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_10_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_10_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_10_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_10_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_10_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_10_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_10_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_10_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_10_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_10_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_in_read : OUT STD_LOGIC;
                    signal nios2_clock_10_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_10_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_10_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_10_in_write : OUT STD_LOGIC;
                    signal nios2_clock_10_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios2_clock_10_in_arbitrator;

component nios2_clock_10_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_mode_select_s1_end_xfer : IN STD_LOGIC;
                    signal mode_select_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_out_granted_mode_select_s1 : IN STD_LOGIC;
                    signal nios2_clock_10_out_qualified_request_mode_select_s1 : IN STD_LOGIC;
                    signal nios2_clock_10_out_read : IN STD_LOGIC;
                    signal nios2_clock_10_out_read_data_valid_mode_select_s1 : IN STD_LOGIC;
                    signal nios2_clock_10_out_requests_mode_select_s1 : IN STD_LOGIC;
                    signal nios2_clock_10_out_write : IN STD_LOGIC;
                    signal nios2_clock_10_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_10_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_10_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_10_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_10_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_10_out_arbitrator;

component nios2_clock_10 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_10;

component nios2_clock_11_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_11_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_11_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_11_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_11_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_11_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_11_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_11_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_11_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_11_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_11_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_11_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_11_in_read : OUT STD_LOGIC;
                    signal nios2_clock_11_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_11_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_11_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_11_in_write : OUT STD_LOGIC;
                    signal nios2_clock_11_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios2_clock_11_in_arbitrator;

component nios2_clock_11_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal comparator_pio_s1_readdata_from_sa : IN STD_LOGIC;
                    signal d1_comparator_pio_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_11_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_11_out_granted_comparator_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_11_out_qualified_request_comparator_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_11_out_read : IN STD_LOGIC;
                    signal nios2_clock_11_out_read_data_valid_comparator_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_11_out_requests_comparator_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_11_out_write : IN STD_LOGIC;
                    signal nios2_clock_11_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_11_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_11_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_11_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_11_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_11_out_arbitrator;

component nios2_clock_11 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_11;

component nios2_clock_12_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_12_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_12_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_12_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_12_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_12_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_12_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_12_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_12_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_12_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_12_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_12_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_12_in_read : OUT STD_LOGIC;
                    signal nios2_clock_12_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_12_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_12_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_12_in_write : OUT STD_LOGIC;
                    signal nios2_clock_12_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios2_clock_12_in_arbitrator;

component nios2_clock_12_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_12_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_12_out_granted_led_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_12_out_qualified_request_led_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_12_out_read : IN STD_LOGIC;
                    signal nios2_clock_12_out_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_12_out_requests_led_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_12_out_write : IN STD_LOGIC;
                    signal nios2_clock_12_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_12_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_12_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_12_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_12_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_12_out_arbitrator;

component nios2_clock_12 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_12;

component nios2_clock_13_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_13_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_13_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_13_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_13_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_13_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_13_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_13_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_13_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_13_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_13_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_13_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_13_in_read : OUT STD_LOGIC;
                    signal nios2_clock_13_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_13_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_13_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_13_in_write : OUT STD_LOGIC;
                    signal nios2_clock_13_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios2_clock_13_in_arbitrator;

component nios2_clock_13_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_gen_code_strobe_s1_end_xfer : IN STD_LOGIC;
                    signal gen_code_strobe_s1_readdata_from_sa : IN STD_LOGIC;
                    signal nios2_clock_13_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_13_out_granted_gen_code_strobe_s1 : IN STD_LOGIC;
                    signal nios2_clock_13_out_qualified_request_gen_code_strobe_s1 : IN STD_LOGIC;
                    signal nios2_clock_13_out_read : IN STD_LOGIC;
                    signal nios2_clock_13_out_read_data_valid_gen_code_strobe_s1 : IN STD_LOGIC;
                    signal nios2_clock_13_out_requests_gen_code_strobe_s1 : IN STD_LOGIC;
                    signal nios2_clock_13_out_write : IN STD_LOGIC;
                    signal nios2_clock_13_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_13_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_13_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_13_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_13_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_13_out_arbitrator;

component nios2_clock_13 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_13;

component nios2_clock_14_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_14_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_14_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_14_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_14_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_14_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_14_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_14_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_14_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_14_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_14_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_14_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_14_in_read : OUT STD_LOGIC;
                    signal nios2_clock_14_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_14_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_14_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_14_in_write : OUT STD_LOGIC;
                    signal nios2_clock_14_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios2_clock_14_in_arbitrator;

component nios2_clock_14_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_switch_pio_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_14_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_14_out_granted_switch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_14_out_qualified_request_switch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_14_out_read : IN STD_LOGIC;
                    signal nios2_clock_14_out_read_data_valid_switch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_14_out_requests_switch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_14_out_write : IN STD_LOGIC;
                    signal nios2_clock_14_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal switch_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal nios2_clock_14_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_14_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_14_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_14_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_14_out_arbitrator;

component nios2_clock_14 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_14;

component nios2_clock_15_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_15_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_15_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_15_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_15_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_15_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_15_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_15_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_15_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_15_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_15_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_15_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_15_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_15_in_read : OUT STD_LOGIC;
                    signal nios2_clock_15_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_15_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_15_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_15_in_write : OUT STD_LOGIC;
                    signal nios2_clock_15_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component nios2_clock_15_in_arbitrator;

component nios2_clock_15_out_arbitrator is 
           port (
                 -- inputs:
                    signal cal_dac_code_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_cal_dac_code_pio_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_15_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_15_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_15_out_granted_cal_dac_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_15_out_read : IN STD_LOGIC;
                    signal nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_15_out_requests_cal_dac_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_15_out_write : IN STD_LOGIC;
                    signal nios2_clock_15_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_15_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_15_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_15_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_15_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_15_out_arbitrator;

component nios2_clock_15 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_15;

component nios2_clock_16_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_16_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_16_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_16_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_16_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_16_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_16_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_16_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_16_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_16_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_16_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_16_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_16_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_16_in_read : OUT STD_LOGIC;
                    signal nios2_clock_16_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_16_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_16_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_16_in_write : OUT STD_LOGIC;
                    signal nios2_clock_16_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_clock_16_in_arbitrator;

component nios2_clock_16_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_usb_code_pio_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_16_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_16_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_16_out_granted_usb_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_16_out_qualified_request_usb_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_16_out_read : IN STD_LOGIC;
                    signal nios2_clock_16_out_read_data_valid_usb_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_16_out_requests_usb_code_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_16_out_write : IN STD_LOGIC;
                    signal nios2_clock_16_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal usb_code_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (20 DOWNTO 0);

                 -- outputs:
                    signal nios2_clock_16_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_16_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_16_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_16_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_16_out_arbitrator;

component nios2_clock_16 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_16;

component nios2_clock_17_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_17_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_17_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_17_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_17_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_17_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_17_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_17_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_17_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_17_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_17_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_17_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_17_in_read : OUT STD_LOGIC;
                    signal nios2_clock_17_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_17_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_17_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_17_in_write : OUT STD_LOGIC;
                    signal nios2_clock_17_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios2_clock_17_in_arbitrator;

component nios2_clock_17_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sample_and_hold_pio_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_17_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_17_out_granted_sample_and_hold_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_17_out_read : IN STD_LOGIC;
                    signal nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_17_out_requests_sample_and_hold_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_17_out_write : IN STD_LOGIC;
                    signal nios2_clock_17_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sample_and_hold_pio_s1_readdata_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_17_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_17_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_17_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_17_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_17_out_arbitrator;

component nios2_clock_17 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_17;

component nios2_clock_18_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_18_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_18_in_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_18_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_18_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_18_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_18_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_18_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_18_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_18_in_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_18_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_18_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_18_in_read : OUT STD_LOGIC;
                    signal nios2_clock_18_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_18_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_18_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_18_in_write : OUT STD_LOGIC;
                    signal nios2_clock_18_in_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component nios2_clock_18_in_arbitrator;

component nios2_clock_18_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_latch_pio_s1_end_xfer : IN STD_LOGIC;
                    signal latch_pio_s1_readdata_from_sa : IN STD_LOGIC;
                    signal nios2_clock_18_out_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_18_out_granted_latch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_18_out_qualified_request_latch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_18_out_read : IN STD_LOGIC;
                    signal nios2_clock_18_out_read_data_valid_latch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_18_out_requests_latch_pio_s1 : IN STD_LOGIC;
                    signal nios2_clock_18_out_write : IN STD_LOGIC;
                    signal nios2_clock_18_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_18_out_address_to_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_18_out_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_clock_18_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_18_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_18_out_arbitrator;

component nios2_clock_18 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_18;

component nios2_clock_2_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_2_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_2_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_2_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_2_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_2_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_2_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_2_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_2_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_2_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_2_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_2_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_2_in_nativeaddress : OUT STD_LOGIC;
                    signal nios2_clock_2_in_read : OUT STD_LOGIC;
                    signal nios2_clock_2_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_2_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_2_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_2_in_write : OUT STD_LOGIC;
                    signal nios2_clock_2_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_clock_2_in_arbitrator;

component nios2_clock_2_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_clock_2_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal nios2_clock_2_out_read : IN STD_LOGIC;
                    signal nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal nios2_clock_2_out_write : IN STD_LOGIC;
                    signal nios2_clock_2_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_2_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_2_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_2_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_2_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_2_out_arbitrator;

component nios2_clock_2 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC;
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC;
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_2;

component nios2_clock_3_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_3_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_3_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_3_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_3_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_3_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_3_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_3_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_3_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_3_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_3_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_3_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_3_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_3_in_read : OUT STD_LOGIC;
                    signal nios2_clock_3_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_3_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_3_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_3_in_write : OUT STD_LOGIC;
                    signal nios2_clock_3_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component nios2_clock_3_in_arbitrator;

component nios2_clock_3_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_3_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_3_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_3_out_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal nios2_clock_3_out_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal nios2_clock_3_out_read : IN STD_LOGIC;
                    signal nios2_clock_3_out_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal nios2_clock_3_out_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal nios2_clock_3_out_write : IN STD_LOGIC;
                    signal nios2_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal nios2_clock_3_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_3_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_3_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_3_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_3_out_arbitrator;

component nios2_clock_3 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_3;

component nios2_clock_4_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_4_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_4_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_4_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_4_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_4_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_4_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_4_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_4_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_4_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_4_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_4_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_4_in_nativeaddress : OUT STD_LOGIC;
                    signal nios2_clock_4_in_read : OUT STD_LOGIC;
                    signal nios2_clock_4_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_4_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_4_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_4_in_write : OUT STD_LOGIC;
                    signal nios2_clock_4_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_clock_4_in_arbitrator;

component nios2_clock_4_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_4_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_4_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_4_out_granted_sysid_control_slave : IN STD_LOGIC;
                    signal nios2_clock_4_out_qualified_request_sysid_control_slave : IN STD_LOGIC;
                    signal nios2_clock_4_out_read : IN STD_LOGIC;
                    signal nios2_clock_4_out_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                    signal nios2_clock_4_out_requests_sysid_control_slave : IN STD_LOGIC;
                    signal nios2_clock_4_out_write : IN STD_LOGIC;
                    signal nios2_clock_4_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal nios2_clock_4_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_4_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_4_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_4_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_4_out_arbitrator;

component nios2_clock_4 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC;
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC;
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_4;

component nios2_clock_5_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_5_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_5_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_5_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_5_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_5_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_5_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_5_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_5_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_5_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_5_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_5_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_5_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_5_in_read : OUT STD_LOGIC;
                    signal nios2_clock_5_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_5_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_5_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_5_in_write : OUT STD_LOGIC;
                    signal nios2_clock_5_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_clock_5_in_arbitrator;

component nios2_clock_5_out_arbitrator is 
           port (
                 -- inputs:
                    signal altpll_0_pll_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_altpll_0_pll_slave_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_5_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_5_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_5_out_granted_altpll_0_pll_slave : IN STD_LOGIC;
                    signal nios2_clock_5_out_qualified_request_altpll_0_pll_slave : IN STD_LOGIC;
                    signal nios2_clock_5_out_read : IN STD_LOGIC;
                    signal nios2_clock_5_out_read_data_valid_altpll_0_pll_slave : IN STD_LOGIC;
                    signal nios2_clock_5_out_requests_altpll_0_pll_slave : IN STD_LOGIC;
                    signal nios2_clock_5_out_write : IN STD_LOGIC;
                    signal nios2_clock_5_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_5_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_5_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_5_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_5_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_5_out_arbitrator;

component nios2_clock_5 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_5;

component nios2_clock_6_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_6_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_6_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_6_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_6_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_6_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_6_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_6_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_6_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_6_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_6_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_6_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_6_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_6_in_read : OUT STD_LOGIC;
                    signal nios2_clock_6_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_6_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_6_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_6_in_write : OUT STD_LOGIC;
                    signal nios2_clock_6_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_clock_6_in_arbitrator;

component nios2_clock_6_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_gen_code_value_pio_0_s1_end_xfer : IN STD_LOGIC;
                    signal gen_code_value_pio_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal nios2_clock_6_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_6_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_6_out_granted_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_6_out_read : IN STD_LOGIC;
                    signal nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_6_out_requests_gen_code_value_pio_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_6_out_write : IN STD_LOGIC;
                    signal nios2_clock_6_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_6_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_6_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_6_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_6_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_6_out_arbitrator;

component nios2_clock_6 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_6;

component nios2_clock_7_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_7_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_7_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_7_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_nios2_clock_7_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_7_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_7_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_7_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_7_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_7_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_7_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_7_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_7_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_7_in_read : OUT STD_LOGIC;
                    signal nios2_clock_7_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_7_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_7_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_7_in_write : OUT STD_LOGIC;
                    signal nios2_clock_7_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_clock_7_in_arbitrator;

component nios2_clock_7_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_gen_code_value_pio_1_s1_end_xfer : IN STD_LOGIC;
                    signal gen_code_value_pio_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal nios2_clock_7_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_7_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_7_out_granted_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                    signal nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                    signal nios2_clock_7_out_read : IN STD_LOGIC;
                    signal nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                    signal nios2_clock_7_out_requests_gen_code_value_pio_1_s1 : IN STD_LOGIC;
                    signal nios2_clock_7_out_write : IN STD_LOGIC;
                    signal nios2_clock_7_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_7_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_7_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_7_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_7_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_7_out_arbitrator;

component nios2_clock_7 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_7;

component nios2_clock_8_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_0_instruction_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal nios2_clock_8_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_8_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_8_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_instruction_master_granted_nios2_clock_8_in : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_nios2_clock_8_in : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_nios2_clock_8_in : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_nios2_clock_8_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_8_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_8_in_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_8_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_8_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_8_in_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal nios2_clock_8_in_read : OUT STD_LOGIC;
                    signal nios2_clock_8_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_8_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_8_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_8_in_write : OUT STD_LOGIC
                 );
end component nios2_clock_8_in_arbitrator;

component nios2_clock_8_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_8_out_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_8_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_8_out_granted_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_8_out_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_8_out_read : IN STD_LOGIC;
                    signal nios2_clock_8_out_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal nios2_clock_8_out_requests_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_8_out_write : IN STD_LOGIC;
                    signal nios2_clock_8_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_8_out_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_8_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_8_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_8_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_8_out_arbitrator;

component nios2_clock_8 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_8;

component nios2_clock_9_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_0_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_0_data_master_latency_counter : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal nios2_clock_9_in_endofpacket : IN STD_LOGIC;
                    signal nios2_clock_9_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_9_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_byteenable_nios2_clock_9_in : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_0_data_master_granted_nios2_clock_9_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_nios2_clock_9_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_nios2_clock_9_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_nios2_clock_9_in : OUT STD_LOGIC;
                    signal d1_nios2_clock_9_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_9_in_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_9_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_9_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_9_in_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal nios2_clock_9_in_read : OUT STD_LOGIC;
                    signal nios2_clock_9_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_9_in_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_9_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_clock_9_in_write : OUT STD_LOGIC;
                    signal nios2_clock_9_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component nios2_clock_9_in_arbitrator;

component nios2_clock_9_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_clock_9_out_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_9_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_9_out_granted_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_9_out_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_9_out_read : IN STD_LOGIC;
                    signal nios2_clock_9_out_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal nios2_clock_9_out_requests_sdram_0_s1 : IN STD_LOGIC;
                    signal nios2_clock_9_out_write : IN STD_LOGIC;
                    signal nios2_clock_9_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_clock_9_out_address_to_slave : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_9_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_9_out_reset_n : OUT STD_LOGIC;
                    signal nios2_clock_9_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_9_out_arbitrator;

component nios2_clock_9 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_clock_9;

component onchip_mem_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_0_out_read : IN STD_LOGIC;
                    signal nios2_clock_0_out_write : IN STD_LOGIC;
                    signal nios2_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_1_out_read : IN STD_LOGIC;
                    signal nios2_clock_1_out_write : IN STD_LOGIC;
                    signal nios2_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal onchip_mem_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_onchip_mem_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_0_out_granted_onchip_mem_s1 : OUT STD_LOGIC;
                    signal nios2_clock_0_out_qualified_request_onchip_mem_s1 : OUT STD_LOGIC;
                    signal nios2_clock_0_out_read_data_valid_onchip_mem_s1 : OUT STD_LOGIC;
                    signal nios2_clock_0_out_requests_onchip_mem_s1 : OUT STD_LOGIC;
                    signal nios2_clock_1_out_granted_onchip_mem_s1 : OUT STD_LOGIC;
                    signal nios2_clock_1_out_qualified_request_onchip_mem_s1 : OUT STD_LOGIC;
                    signal nios2_clock_1_out_read_data_valid_onchip_mem_s1 : OUT STD_LOGIC;
                    signal nios2_clock_1_out_requests_onchip_mem_s1 : OUT STD_LOGIC;
                    signal onchip_mem_s1_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal onchip_mem_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal onchip_mem_s1_chipselect : OUT STD_LOGIC;
                    signal onchip_mem_s1_clken : OUT STD_LOGIC;
                    signal onchip_mem_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal onchip_mem_s1_reset : OUT STD_LOGIC;
                    signal onchip_mem_s1_write : OUT STD_LOGIC;
                    signal onchip_mem_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component onchip_mem_s1_arbitrator;

component onchip_mem is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component onchip_mem;

component sample_and_hold_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_17_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_17_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_17_out_read : IN STD_LOGIC;
                    signal nios2_clock_17_out_write : IN STD_LOGIC;
                    signal nios2_clock_17_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sample_and_hold_pio_s1_readdata : IN STD_LOGIC;

                 -- outputs:
                    signal d1_sample_and_hold_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_17_out_granted_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_17_out_requests_sample_and_hold_pio_s1 : OUT STD_LOGIC;
                    signal sample_and_hold_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sample_and_hold_pio_s1_chipselect : OUT STD_LOGIC;
                    signal sample_and_hold_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal sample_and_hold_pio_s1_reset_n : OUT STD_LOGIC;
                    signal sample_and_hold_pio_s1_write_n : OUT STD_LOGIC;
                    signal sample_and_hold_pio_s1_writedata : OUT STD_LOGIC
                 );
end component sample_and_hold_pio_s1_arbitrator;

component sample_and_hold_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component sample_and_hold_pio;

component sdram_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_8_out_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_8_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_8_out_read : IN STD_LOGIC;
                    signal nios2_clock_8_out_write : IN STD_LOGIC;
                    signal nios2_clock_8_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_clock_9_out_address_to_slave : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal nios2_clock_9_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_9_out_read : IN STD_LOGIC;
                    signal nios2_clock_9_out_write : IN STD_LOGIC;
                    signal nios2_clock_9_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_0_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_0_s1_readdatavalid : IN STD_LOGIC;
                    signal sdram_0_s1_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal d1_sdram_0_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_8_out_granted_sdram_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_8_out_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_8_out_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                    signal nios2_clock_8_out_requests_sdram_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_9_out_granted_sdram_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_9_out_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_9_out_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                    signal nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                    signal nios2_clock_9_out_requests_sdram_0_s1 : OUT STD_LOGIC;
                    signal sdram_0_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal sdram_0_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sdram_0_s1_chipselect : OUT STD_LOGIC;
                    signal sdram_0_s1_read_n : OUT STD_LOGIC;
                    signal sdram_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_0_s1_reset_n : OUT STD_LOGIC;
                    signal sdram_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal sdram_0_s1_write_n : OUT STD_LOGIC;
                    signal sdram_0_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sdram_0_s1_arbitrator;

component sdram_0 is 
           port (
                 -- inputs:
                    signal az_addr : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal az_be_n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal az_cs : IN STD_LOGIC;
                    signal az_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal az_rd_n : IN STD_LOGIC;
                    signal az_wr_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal za_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal za_valid : OUT STD_LOGIC;
                    signal za_waitrequest : OUT STD_LOGIC;
                    signal zs_addr : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : OUT STD_LOGIC;
                    signal zs_cke : OUT STD_LOGIC;
                    signal zs_cs_n : OUT STD_LOGIC;
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n : OUT STD_LOGIC;
                    signal zs_we_n : OUT STD_LOGIC
                 );
end component sdram_0;

component switch_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_14_out_address_to_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_14_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_14_out_read : IN STD_LOGIC;
                    signal nios2_clock_14_out_write : IN STD_LOGIC;
                    signal nios2_clock_14_out_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal switch_pio_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal d1_switch_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_14_out_granted_switch_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_14_out_qualified_request_switch_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_14_out_read_data_valid_switch_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_14_out_requests_switch_pio_s1 : OUT STD_LOGIC;
                    signal switch_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal switch_pio_s1_chipselect : OUT STD_LOGIC;
                    signal switch_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal switch_pio_s1_reset_n : OUT STD_LOGIC;
                    signal switch_pio_s1_write_n : OUT STD_LOGIC;
                    signal switch_pio_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component switch_pio_s1_arbitrator;

component switch_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component switch_pio;

component sys_clk_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_3_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_3_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_3_out_read : IN STD_LOGIC;
                    signal nios2_clock_3_out_write : IN STD_LOGIC;
                    signal nios2_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                    signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_3_out_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal nios2_clock_3_out_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal nios2_clock_3_out_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal nios2_clock_3_out_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer_s1_arbitrator;

component sys_clk_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer;

component sysid_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_4_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_clock_4_out_nativeaddress : IN STD_LOGIC;
                    signal nios2_clock_4_out_read : IN STD_LOGIC;
                    signal nios2_clock_4_out_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_4_out_granted_sysid_control_slave : OUT STD_LOGIC;
                    signal nios2_clock_4_out_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                    signal nios2_clock_4_out_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                    signal nios2_clock_4_out_requests_sysid_control_slave : OUT STD_LOGIC;
                    signal sysid_control_slave_address : OUT STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sysid_control_slave_reset_n : OUT STD_LOGIC
                 );
end component sysid_control_slave_arbitrator;

component sysid is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;
                    signal clock : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid;

component usb_code_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_clock_16_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_clock_16_out_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_clock_16_out_read : IN STD_LOGIC;
                    signal nios2_clock_16_out_write : IN STD_LOGIC;
                    signal nios2_clock_16_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal usb_code_pio_s1_readdata : IN STD_LOGIC_VECTOR (20 DOWNTO 0);

                 -- outputs:
                    signal d1_usb_code_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_clock_16_out_granted_usb_code_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_16_out_qualified_request_usb_code_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_16_out_read_data_valid_usb_code_pio_s1 : OUT STD_LOGIC;
                    signal nios2_clock_16_out_requests_usb_code_pio_s1 : OUT STD_LOGIC;
                    signal usb_code_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal usb_code_pio_s1_chipselect : OUT STD_LOGIC;
                    signal usb_code_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal usb_code_pio_s1_reset_n : OUT STD_LOGIC;
                    signal usb_code_pio_s1_write_n : OUT STD_LOGIC;
                    signal usb_code_pio_s1_writedata : OUT STD_LOGIC_VECTOR (20 DOWNTO 0)
                 );
end component usb_code_pio_s1_arbitrator;

component usb_code_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (20 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (20 DOWNTO 0)
                 );
end component usb_code_pio;

component nios2_reset_clk_0_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios2_reset_clk_0_domain_synch_module;

component nios2_reset_altpll_0_c0_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios2_reset_altpll_0_c0_domain_synch_module;

component nios2_reset_processor_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios2_reset_processor_clk_domain_synch_module;

component nios2_reset_altpll_0_c1_out_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios2_reset_altpll_0_c1_out_domain_synch_module;

                signal altpll_0_c0_reset_n :  STD_LOGIC;
                signal altpll_0_c1_out_reset_n :  STD_LOGIC;
                signal altpll_0_pll_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal altpll_0_pll_slave_read :  STD_LOGIC;
                signal altpll_0_pll_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal altpll_0_pll_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal altpll_0_pll_slave_reset :  STD_LOGIC;
                signal altpll_0_pll_slave_write :  STD_LOGIC;
                signal altpll_0_pll_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cal_dac_code_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cal_dac_code_pio_s1_chipselect :  STD_LOGIC;
                signal cal_dac_code_pio_s1_readdata :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal cal_dac_code_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal cal_dac_code_pio_s1_reset_n :  STD_LOGIC;
                signal cal_dac_code_pio_s1_write_n :  STD_LOGIC;
                signal cal_dac_code_pio_s1_writedata :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal clk_0_reset_n :  STD_LOGIC;
                signal comparator_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal comparator_pio_s1_readdata :  STD_LOGIC;
                signal comparator_pio_s1_readdata_from_sa :  STD_LOGIC;
                signal comparator_pio_s1_reset_n :  STD_LOGIC;
                signal cpu_0_data_master_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_0_data_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_0_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_0_data_master_byteenable_nios2_clock_9_in :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_data_master_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal cpu_0_data_master_debugaccess :  STD_LOGIC;
                signal cpu_0_data_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_10_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_11_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_12_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_13_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_14_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_15_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_16_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_17_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_18_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_2_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_3_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_4_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_5_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_6_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_7_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_nios2_clock_9_in :  STD_LOGIC;
                signal cpu_0_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_data_master_latency_counter :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_10_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_11_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_12_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_13_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_14_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_15_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_16_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_17_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_18_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_2_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_3_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_4_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_5_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_6_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_7_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_nios2_clock_9_in :  STD_LOGIC;
                signal cpu_0_data_master_read :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_10_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_11_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_12_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_13_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_14_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_15_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_16_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_17_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_18_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_2_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_3_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_4_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_5_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_6_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_7_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_nios2_clock_9_in :  STD_LOGIC;
                signal cpu_0_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_data_master_readdatavalid :  STD_LOGIC;
                signal cpu_0_data_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_10_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_11_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_12_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_13_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_14_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_15_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_16_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_17_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_18_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_2_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_3_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_4_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_5_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_6_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_7_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_nios2_clock_9_in :  STD_LOGIC;
                signal cpu_0_data_master_waitrequest :  STD_LOGIC;
                signal cpu_0_data_master_write :  STD_LOGIC;
                signal cpu_0_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_instruction_master_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_0_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_0_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_granted_nios2_clock_0_in :  STD_LOGIC;
                signal cpu_0_instruction_master_granted_nios2_clock_8_in :  STD_LOGIC;
                signal cpu_0_instruction_master_latency_counter :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_nios2_clock_0_in :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_nios2_clock_8_in :  STD_LOGIC;
                signal cpu_0_instruction_master_read :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_nios2_clock_0_in :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_nios2_clock_8_in :  STD_LOGIC;
                signal cpu_0_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_instruction_master_readdatavalid :  STD_LOGIC;
                signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_requests_nios2_clock_0_in :  STD_LOGIC;
                signal cpu_0_instruction_master_requests_nios2_clock_8_in :  STD_LOGIC;
                signal cpu_0_instruction_master_waitrequest :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal cpu_0_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_0_jtag_debug_module_chipselect :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_jtag_debug_module_reset_n :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_write :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_altpll_0_pll_slave_end_xfer :  STD_LOGIC;
                signal d1_cal_dac_code_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_comparator_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_cpu_0_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_gen_code_strobe_s1_end_xfer :  STD_LOGIC;
                signal d1_gen_code_value_pio_0_s1_end_xfer :  STD_LOGIC;
                signal d1_gen_code_value_pio_1_s1_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_latch_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_led_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_mode_select_s1_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_0_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_10_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_11_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_12_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_13_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_14_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_15_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_16_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_17_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_18_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_1_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_2_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_3_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_4_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_5_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_6_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_7_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_8_in_end_xfer :  STD_LOGIC;
                signal d1_nios2_clock_9_in_end_xfer :  STD_LOGIC;
                signal d1_onchip_mem_s1_end_xfer :  STD_LOGIC;
                signal d1_sample_and_hold_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_sdram_0_s1_end_xfer :  STD_LOGIC;
                signal d1_switch_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_sysid_control_slave_end_xfer :  STD_LOGIC;
                signal d1_usb_code_pio_s1_end_xfer :  STD_LOGIC;
                signal gen_code_strobe_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gen_code_strobe_s1_chipselect :  STD_LOGIC;
                signal gen_code_strobe_s1_readdata :  STD_LOGIC;
                signal gen_code_strobe_s1_readdata_from_sa :  STD_LOGIC;
                signal gen_code_strobe_s1_reset_n :  STD_LOGIC;
                signal gen_code_strobe_s1_write_n :  STD_LOGIC;
                signal gen_code_strobe_s1_writedata :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gen_code_value_pio_0_s1_chipselect :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_readdata :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal gen_code_value_pio_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal gen_code_value_pio_0_s1_reset_n :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_write_n :  STD_LOGIC;
                signal gen_code_value_pio_0_s1_writedata :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal gen_code_value_pio_1_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gen_code_value_pio_1_s1_chipselect :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_readdata :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal gen_code_value_pio_1_s1_readdata_from_sa :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal gen_code_value_pio_1_s1_reset_n :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_write_n :  STD_LOGIC;
                signal gen_code_value_pio_1_s1_writedata :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal internal_altpll_0_c0 :  STD_LOGIC;
                signal internal_altpll_0_c1_out :  STD_LOGIC;
                signal internal_locked_from_the_altpll_0 :  STD_LOGIC;
                signal internal_out_port_from_the_cal_dac_code_pio :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal internal_out_port_from_the_gen_code_strobe :  STD_LOGIC;
                signal internal_out_port_from_the_gen_code_value_pio_0 :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal internal_out_port_from_the_gen_code_value_pio_1 :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal internal_out_port_from_the_latch_pio :  STD_LOGIC;
                signal internal_out_port_from_the_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_sample_and_hold_pio :  STD_LOGIC;
                signal internal_out_port_from_the_switch_pio :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_out_port_from_the_usb_code_pio :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal internal_phasedone_from_the_altpll_0 :  STD_LOGIC;
                signal internal_zs_addr_from_the_sdram_0 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal internal_zs_ba_from_the_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_cas_n_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_cke_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_cs_n_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_dqm_from_the_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_ras_n_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_we_n_from_the_sdram_0 :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_0_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal latch_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal latch_pio_s1_chipselect :  STD_LOGIC;
                signal latch_pio_s1_readdata :  STD_LOGIC;
                signal latch_pio_s1_readdata_from_sa :  STD_LOGIC;
                signal latch_pio_s1_reset_n :  STD_LOGIC;
                signal latch_pio_s1_write_n :  STD_LOGIC;
                signal latch_pio_s1_writedata :  STD_LOGIC;
                signal led_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal led_pio_s1_chipselect :  STD_LOGIC;
                signal led_pio_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_reset_n :  STD_LOGIC;
                signal led_pio_s1_write_n :  STD_LOGIC;
                signal led_pio_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal mode_select_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mode_select_s1_chipselect :  STD_LOGIC;
                signal mode_select_s1_readdata :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mode_select_s1_readdata_from_sa :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mode_select_s1_reset_n :  STD_LOGIC;
                signal mode_select_s1_write_n :  STD_LOGIC;
                signal mode_select_s1_writedata :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal nios2_clock_0_in_address :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_0_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_0_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_0_in_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_clock_0_in_read :  STD_LOGIC;
                signal nios2_clock_0_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_0_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_0_in_reset_n :  STD_LOGIC;
                signal nios2_clock_0_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_0_in_write :  STD_LOGIC;
                signal nios2_clock_0_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_0_out_address :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_0_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_0_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_0_out_granted_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_0_out_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_clock_0_out_qualified_request_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_0_out_read :  STD_LOGIC;
                signal nios2_clock_0_out_read_data_valid_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_0_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_0_out_requests_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_0_out_reset_n :  STD_LOGIC;
                signal nios2_clock_0_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_0_out_write :  STD_LOGIC;
                signal nios2_clock_0_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_10_in_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_10_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_10_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_in_read :  STD_LOGIC;
                signal nios2_clock_10_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_10_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_10_in_reset_n :  STD_LOGIC;
                signal nios2_clock_10_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_10_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_10_in_write :  STD_LOGIC;
                signal nios2_clock_10_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_10_out_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_10_out_granted_mode_select_s1 :  STD_LOGIC;
                signal nios2_clock_10_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_10_out_qualified_request_mode_select_s1 :  STD_LOGIC;
                signal nios2_clock_10_out_read :  STD_LOGIC;
                signal nios2_clock_10_out_read_data_valid_mode_select_s1 :  STD_LOGIC;
                signal nios2_clock_10_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_10_out_requests_mode_select_s1 :  STD_LOGIC;
                signal nios2_clock_10_out_reset_n :  STD_LOGIC;
                signal nios2_clock_10_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_10_out_write :  STD_LOGIC;
                signal nios2_clock_10_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_11_in_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_11_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_11_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_in_read :  STD_LOGIC;
                signal nios2_clock_11_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_11_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_11_in_reset_n :  STD_LOGIC;
                signal nios2_clock_11_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_11_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_11_in_write :  STD_LOGIC;
                signal nios2_clock_11_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_11_out_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_11_out_granted_comparator_pio_s1 :  STD_LOGIC;
                signal nios2_clock_11_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_11_out_qualified_request_comparator_pio_s1 :  STD_LOGIC;
                signal nios2_clock_11_out_read :  STD_LOGIC;
                signal nios2_clock_11_out_read_data_valid_comparator_pio_s1 :  STD_LOGIC;
                signal nios2_clock_11_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_11_out_requests_comparator_pio_s1 :  STD_LOGIC;
                signal nios2_clock_11_out_reset_n :  STD_LOGIC;
                signal nios2_clock_11_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_11_out_write :  STD_LOGIC;
                signal nios2_clock_11_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_12_in_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_12_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_12_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_in_read :  STD_LOGIC;
                signal nios2_clock_12_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_12_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_12_in_reset_n :  STD_LOGIC;
                signal nios2_clock_12_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_12_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_12_in_write :  STD_LOGIC;
                signal nios2_clock_12_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_12_out_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_12_out_granted_led_pio_s1 :  STD_LOGIC;
                signal nios2_clock_12_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_12_out_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal nios2_clock_12_out_read :  STD_LOGIC;
                signal nios2_clock_12_out_read_data_valid_led_pio_s1 :  STD_LOGIC;
                signal nios2_clock_12_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_12_out_requests_led_pio_s1 :  STD_LOGIC;
                signal nios2_clock_12_out_reset_n :  STD_LOGIC;
                signal nios2_clock_12_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_12_out_write :  STD_LOGIC;
                signal nios2_clock_12_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_13_in_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_13_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_13_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_in_read :  STD_LOGIC;
                signal nios2_clock_13_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_13_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_13_in_reset_n :  STD_LOGIC;
                signal nios2_clock_13_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_13_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_13_in_write :  STD_LOGIC;
                signal nios2_clock_13_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_13_out_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_13_out_granted_gen_code_strobe_s1 :  STD_LOGIC;
                signal nios2_clock_13_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_13_out_qualified_request_gen_code_strobe_s1 :  STD_LOGIC;
                signal nios2_clock_13_out_read :  STD_LOGIC;
                signal nios2_clock_13_out_read_data_valid_gen_code_strobe_s1 :  STD_LOGIC;
                signal nios2_clock_13_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_13_out_requests_gen_code_strobe_s1 :  STD_LOGIC;
                signal nios2_clock_13_out_reset_n :  STD_LOGIC;
                signal nios2_clock_13_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_13_out_write :  STD_LOGIC;
                signal nios2_clock_13_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_14_in_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_14_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_14_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_in_read :  STD_LOGIC;
                signal nios2_clock_14_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_14_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_14_in_reset_n :  STD_LOGIC;
                signal nios2_clock_14_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_14_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_14_in_write :  STD_LOGIC;
                signal nios2_clock_14_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_14_out_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_14_out_granted_switch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_14_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_14_out_qualified_request_switch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_14_out_read :  STD_LOGIC;
                signal nios2_clock_14_out_read_data_valid_switch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_14_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_14_out_requests_switch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_14_out_reset_n :  STD_LOGIC;
                signal nios2_clock_14_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_14_out_write :  STD_LOGIC;
                signal nios2_clock_14_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_15_in_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_15_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_15_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_15_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_in_read :  STD_LOGIC;
                signal nios2_clock_15_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_15_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_15_in_reset_n :  STD_LOGIC;
                signal nios2_clock_15_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_15_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_15_in_write :  STD_LOGIC;
                signal nios2_clock_15_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_15_out_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_15_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_15_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_15_out_granted_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_15_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_15_out_read :  STD_LOGIC;
                signal nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_15_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_15_out_requests_cal_dac_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_15_out_reset_n :  STD_LOGIC;
                signal nios2_clock_15_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_15_out_write :  STD_LOGIC;
                signal nios2_clock_15_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_16_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_16_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_16_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_16_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_16_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_16_in_read :  STD_LOGIC;
                signal nios2_clock_16_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_16_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_16_in_reset_n :  STD_LOGIC;
                signal nios2_clock_16_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_16_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_16_in_write :  STD_LOGIC;
                signal nios2_clock_16_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_16_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_16_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_16_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_16_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_16_out_granted_usb_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_16_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_16_out_qualified_request_usb_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_16_out_read :  STD_LOGIC;
                signal nios2_clock_16_out_read_data_valid_usb_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_16_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_16_out_requests_usb_code_pio_s1 :  STD_LOGIC;
                signal nios2_clock_16_out_reset_n :  STD_LOGIC;
                signal nios2_clock_16_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_16_out_write :  STD_LOGIC;
                signal nios2_clock_16_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_17_in_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_17_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_17_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_in_read :  STD_LOGIC;
                signal nios2_clock_17_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_17_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_17_in_reset_n :  STD_LOGIC;
                signal nios2_clock_17_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_17_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_17_in_write :  STD_LOGIC;
                signal nios2_clock_17_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_17_out_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_17_out_granted_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal nios2_clock_17_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal nios2_clock_17_out_read :  STD_LOGIC;
                signal nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal nios2_clock_17_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_17_out_requests_sample_and_hold_pio_s1 :  STD_LOGIC;
                signal nios2_clock_17_out_reset_n :  STD_LOGIC;
                signal nios2_clock_17_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_17_out_write :  STD_LOGIC;
                signal nios2_clock_17_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_18_in_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_18_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_18_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_in_read :  STD_LOGIC;
                signal nios2_clock_18_in_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_18_in_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_18_in_reset_n :  STD_LOGIC;
                signal nios2_clock_18_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_18_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_18_in_write :  STD_LOGIC;
                signal nios2_clock_18_in_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_18_out_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_out_address_to_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_18_out_granted_latch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_18_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_18_out_qualified_request_latch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_18_out_read :  STD_LOGIC;
                signal nios2_clock_18_out_read_data_valid_latch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_18_out_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_18_out_requests_latch_pio_s1 :  STD_LOGIC;
                signal nios2_clock_18_out_reset_n :  STD_LOGIC;
                signal nios2_clock_18_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_18_out_write :  STD_LOGIC;
                signal nios2_clock_18_out_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_clock_1_in_address :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_1_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_1_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_1_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_1_in_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_clock_1_in_read :  STD_LOGIC;
                signal nios2_clock_1_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_1_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_1_in_reset_n :  STD_LOGIC;
                signal nios2_clock_1_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_1_in_write :  STD_LOGIC;
                signal nios2_clock_1_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_1_out_address :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_clock_1_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_1_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_1_out_granted_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_1_out_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_clock_1_out_qualified_request_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_1_out_read :  STD_LOGIC;
                signal nios2_clock_1_out_read_data_valid_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_1_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_1_out_requests_onchip_mem_s1 :  STD_LOGIC;
                signal nios2_clock_1_out_reset_n :  STD_LOGIC;
                signal nios2_clock_1_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_1_out_write :  STD_LOGIC;
                signal nios2_clock_1_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_2_in_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_2_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_2_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_2_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_2_in_nativeaddress :  STD_LOGIC;
                signal nios2_clock_2_in_read :  STD_LOGIC;
                signal nios2_clock_2_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_2_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_2_in_reset_n :  STD_LOGIC;
                signal nios2_clock_2_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_2_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_2_in_write :  STD_LOGIC;
                signal nios2_clock_2_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_2_out_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_2_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_2_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_2_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal nios2_clock_2_out_nativeaddress :  STD_LOGIC;
                signal nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal nios2_clock_2_out_read :  STD_LOGIC;
                signal nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal nios2_clock_2_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal nios2_clock_2_out_reset_n :  STD_LOGIC;
                signal nios2_clock_2_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_2_out_write :  STD_LOGIC;
                signal nios2_clock_2_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_3_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_3_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_3_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_3_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_3_in_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_3_in_read :  STD_LOGIC;
                signal nios2_clock_3_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_3_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_3_in_reset_n :  STD_LOGIC;
                signal nios2_clock_3_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_3_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_3_in_write :  STD_LOGIC;
                signal nios2_clock_3_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_3_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_3_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_3_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_3_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_3_out_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal nios2_clock_3_out_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_3_out_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal nios2_clock_3_out_read :  STD_LOGIC;
                signal nios2_clock_3_out_read_data_valid_sys_clk_timer_s1 :  STD_LOGIC;
                signal nios2_clock_3_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_3_out_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal nios2_clock_3_out_reset_n :  STD_LOGIC;
                signal nios2_clock_3_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_3_out_write :  STD_LOGIC;
                signal nios2_clock_3_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_4_in_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_4_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_4_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_4_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_4_in_nativeaddress :  STD_LOGIC;
                signal nios2_clock_4_in_read :  STD_LOGIC;
                signal nios2_clock_4_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_4_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_4_in_reset_n :  STD_LOGIC;
                signal nios2_clock_4_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_4_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_4_in_write :  STD_LOGIC;
                signal nios2_clock_4_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_4_out_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_4_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_clock_4_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_4_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_4_out_granted_sysid_control_slave :  STD_LOGIC;
                signal nios2_clock_4_out_nativeaddress :  STD_LOGIC;
                signal nios2_clock_4_out_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal nios2_clock_4_out_read :  STD_LOGIC;
                signal nios2_clock_4_out_read_data_valid_sysid_control_slave :  STD_LOGIC;
                signal nios2_clock_4_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_4_out_requests_sysid_control_slave :  STD_LOGIC;
                signal nios2_clock_4_out_reset_n :  STD_LOGIC;
                signal nios2_clock_4_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_4_out_write :  STD_LOGIC;
                signal nios2_clock_4_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_5_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_5_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_5_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_5_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_5_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_5_in_read :  STD_LOGIC;
                signal nios2_clock_5_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_5_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_5_in_reset_n :  STD_LOGIC;
                signal nios2_clock_5_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_5_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_5_in_write :  STD_LOGIC;
                signal nios2_clock_5_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_5_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_5_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_5_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_5_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_5_out_granted_altpll_0_pll_slave :  STD_LOGIC;
                signal nios2_clock_5_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_5_out_qualified_request_altpll_0_pll_slave :  STD_LOGIC;
                signal nios2_clock_5_out_read :  STD_LOGIC;
                signal nios2_clock_5_out_read_data_valid_altpll_0_pll_slave :  STD_LOGIC;
                signal nios2_clock_5_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_5_out_requests_altpll_0_pll_slave :  STD_LOGIC;
                signal nios2_clock_5_out_reset_n :  STD_LOGIC;
                signal nios2_clock_5_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_5_out_write :  STD_LOGIC;
                signal nios2_clock_5_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_6_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_6_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_6_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_6_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_6_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_6_in_read :  STD_LOGIC;
                signal nios2_clock_6_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_6_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_6_in_reset_n :  STD_LOGIC;
                signal nios2_clock_6_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_6_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_6_in_write :  STD_LOGIC;
                signal nios2_clock_6_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_6_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_6_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_6_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_6_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_6_out_granted_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal nios2_clock_6_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal nios2_clock_6_out_read :  STD_LOGIC;
                signal nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal nios2_clock_6_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_6_out_requests_gen_code_value_pio_0_s1 :  STD_LOGIC;
                signal nios2_clock_6_out_reset_n :  STD_LOGIC;
                signal nios2_clock_6_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_6_out_write :  STD_LOGIC;
                signal nios2_clock_6_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_7_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_7_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_7_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_7_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_7_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_7_in_read :  STD_LOGIC;
                signal nios2_clock_7_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_7_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_7_in_reset_n :  STD_LOGIC;
                signal nios2_clock_7_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_7_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_7_in_write :  STD_LOGIC;
                signal nios2_clock_7_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_7_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_7_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_7_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_clock_7_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_7_out_granted_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal nios2_clock_7_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal nios2_clock_7_out_read :  STD_LOGIC;
                signal nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal nios2_clock_7_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_7_out_requests_gen_code_value_pio_1_s1 :  STD_LOGIC;
                signal nios2_clock_7_out_reset_n :  STD_LOGIC;
                signal nios2_clock_7_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_7_out_write :  STD_LOGIC;
                signal nios2_clock_7_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_8_in_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_8_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_8_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_8_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_8_in_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal nios2_clock_8_in_read :  STD_LOGIC;
                signal nios2_clock_8_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_8_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_8_in_reset_n :  STD_LOGIC;
                signal nios2_clock_8_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_8_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_8_in_write :  STD_LOGIC;
                signal nios2_clock_8_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_8_out_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_8_out_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_8_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_8_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_8_out_granted_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_8_out_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal nios2_clock_8_out_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_8_out_read :  STD_LOGIC;
                signal nios2_clock_8_out_read_data_valid_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register :  STD_LOGIC;
                signal nios2_clock_8_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_8_out_requests_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_8_out_reset_n :  STD_LOGIC;
                signal nios2_clock_8_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_8_out_write :  STD_LOGIC;
                signal nios2_clock_8_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_9_in_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_9_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_9_in_endofpacket :  STD_LOGIC;
                signal nios2_clock_9_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_9_in_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal nios2_clock_9_in_read :  STD_LOGIC;
                signal nios2_clock_9_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_9_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_9_in_reset_n :  STD_LOGIC;
                signal nios2_clock_9_in_waitrequest :  STD_LOGIC;
                signal nios2_clock_9_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_clock_9_in_write :  STD_LOGIC;
                signal nios2_clock_9_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_9_out_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_9_out_address_to_slave :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal nios2_clock_9_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_9_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_9_out_granted_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_9_out_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal nios2_clock_9_out_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_9_out_read :  STD_LOGIC;
                signal nios2_clock_9_out_read_data_valid_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register :  STD_LOGIC;
                signal nios2_clock_9_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_9_out_requests_sdram_0_s1 :  STD_LOGIC;
                signal nios2_clock_9_out_reset_n :  STD_LOGIC;
                signal nios2_clock_9_out_waitrequest :  STD_LOGIC;
                signal nios2_clock_9_out_write :  STD_LOGIC;
                signal nios2_clock_9_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal onchip_mem_s1_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal onchip_mem_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal onchip_mem_s1_chipselect :  STD_LOGIC;
                signal onchip_mem_s1_clken :  STD_LOGIC;
                signal onchip_mem_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal onchip_mem_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal onchip_mem_s1_reset :  STD_LOGIC;
                signal onchip_mem_s1_write :  STD_LOGIC;
                signal onchip_mem_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal out_clk_altpll_0_c0 :  STD_LOGIC;
                signal out_clk_altpll_0_c1 :  STD_LOGIC;
                signal processor_clk_reset_n :  STD_LOGIC;
                signal reset_n_sources :  STD_LOGIC;
                signal sample_and_hold_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sample_and_hold_pio_s1_chipselect :  STD_LOGIC;
                signal sample_and_hold_pio_s1_readdata :  STD_LOGIC;
                signal sample_and_hold_pio_s1_readdata_from_sa :  STD_LOGIC;
                signal sample_and_hold_pio_s1_reset_n :  STD_LOGIC;
                signal sample_and_hold_pio_s1_write_n :  STD_LOGIC;
                signal sample_and_hold_pio_s1_writedata :  STD_LOGIC;
                signal sdram_0_s1_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal sdram_0_s1_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_chipselect :  STD_LOGIC;
                signal sdram_0_s1_read_n :  STD_LOGIC;
                signal sdram_0_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_0_s1_readdatavalid :  STD_LOGIC;
                signal sdram_0_s1_reset_n :  STD_LOGIC;
                signal sdram_0_s1_waitrequest :  STD_LOGIC;
                signal sdram_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal sdram_0_s1_write_n :  STD_LOGIC;
                signal sdram_0_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal switch_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal switch_pio_s1_chipselect :  STD_LOGIC;
                signal switch_pio_s1_readdata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal switch_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal switch_pio_s1_reset_n :  STD_LOGIC;
                signal switch_pio_s1_write_n :  STD_LOGIC;
                signal switch_pio_s1_writedata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sys_clk_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_timer_s1_chipselect :  STD_LOGIC;
                signal sys_clk_timer_s1_irq :  STD_LOGIC;
                signal sys_clk_timer_s1_irq_from_sa :  STD_LOGIC;
                signal sys_clk_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_reset_n :  STD_LOGIC;
                signal sys_clk_timer_s1_write_n :  STD_LOGIC;
                signal sys_clk_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sysid_control_slave_address :  STD_LOGIC;
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal sysid_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_reset_n :  STD_LOGIC;
                signal usb_code_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal usb_code_pio_s1_chipselect :  STD_LOGIC;
                signal usb_code_pio_s1_readdata :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal usb_code_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal usb_code_pio_s1_reset_n :  STD_LOGIC;
                signal usb_code_pio_s1_write_n :  STD_LOGIC;
                signal usb_code_pio_s1_writedata :  STD_LOGIC_VECTOR (20 DOWNTO 0);

begin

  --the_altpll_0_pll_slave, which is an e_instance
  the_altpll_0_pll_slave : altpll_0_pll_slave_arbitrator
    port map(
      altpll_0_pll_slave_address => altpll_0_pll_slave_address,
      altpll_0_pll_slave_read => altpll_0_pll_slave_read,
      altpll_0_pll_slave_readdata_from_sa => altpll_0_pll_slave_readdata_from_sa,
      altpll_0_pll_slave_reset => altpll_0_pll_slave_reset,
      altpll_0_pll_slave_write => altpll_0_pll_slave_write,
      altpll_0_pll_slave_writedata => altpll_0_pll_slave_writedata,
      d1_altpll_0_pll_slave_end_xfer => d1_altpll_0_pll_slave_end_xfer,
      nios2_clock_5_out_granted_altpll_0_pll_slave => nios2_clock_5_out_granted_altpll_0_pll_slave,
      nios2_clock_5_out_qualified_request_altpll_0_pll_slave => nios2_clock_5_out_qualified_request_altpll_0_pll_slave,
      nios2_clock_5_out_read_data_valid_altpll_0_pll_slave => nios2_clock_5_out_read_data_valid_altpll_0_pll_slave,
      nios2_clock_5_out_requests_altpll_0_pll_slave => nios2_clock_5_out_requests_altpll_0_pll_slave,
      altpll_0_pll_slave_readdata => altpll_0_pll_slave_readdata,
      clk => clk_0,
      nios2_clock_5_out_address_to_slave => nios2_clock_5_out_address_to_slave,
      nios2_clock_5_out_read => nios2_clock_5_out_read,
      nios2_clock_5_out_write => nios2_clock_5_out_write,
      nios2_clock_5_out_writedata => nios2_clock_5_out_writedata,
      reset_n => clk_0_reset_n
    );


  --altpll_0_c0 out_clk assignment, which is an e_assign
  internal_altpll_0_c0 <= out_clk_altpll_0_c0;
  --altpll_0_c1_out out_clk assignment, which is an e_assign
  internal_altpll_0_c1_out <= out_clk_altpll_0_c1;
  --the_altpll_0, which is an e_ptf_instance
  the_altpll_0 : altpll_0
    port map(
      c0 => out_clk_altpll_0_c0,
      c1 => out_clk_altpll_0_c1,
      locked => internal_locked_from_the_altpll_0,
      phasedone => internal_phasedone_from_the_altpll_0,
      readdata => altpll_0_pll_slave_readdata,
      address => altpll_0_pll_slave_address,
      clk => clk_0,
      read => altpll_0_pll_slave_read,
      reset => altpll_0_pll_slave_reset,
      write => altpll_0_pll_slave_write,
      writedata => altpll_0_pll_slave_writedata
    );


  --the_cal_dac_code_pio_s1, which is an e_instance
  the_cal_dac_code_pio_s1 : cal_dac_code_pio_s1_arbitrator
    port map(
      cal_dac_code_pio_s1_address => cal_dac_code_pio_s1_address,
      cal_dac_code_pio_s1_chipselect => cal_dac_code_pio_s1_chipselect,
      cal_dac_code_pio_s1_readdata_from_sa => cal_dac_code_pio_s1_readdata_from_sa,
      cal_dac_code_pio_s1_reset_n => cal_dac_code_pio_s1_reset_n,
      cal_dac_code_pio_s1_write_n => cal_dac_code_pio_s1_write_n,
      cal_dac_code_pio_s1_writedata => cal_dac_code_pio_s1_writedata,
      d1_cal_dac_code_pio_s1_end_xfer => d1_cal_dac_code_pio_s1_end_xfer,
      nios2_clock_15_out_granted_cal_dac_code_pio_s1 => nios2_clock_15_out_granted_cal_dac_code_pio_s1,
      nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 => nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1,
      nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1 => nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1,
      nios2_clock_15_out_requests_cal_dac_code_pio_s1 => nios2_clock_15_out_requests_cal_dac_code_pio_s1,
      cal_dac_code_pio_s1_readdata => cal_dac_code_pio_s1_readdata,
      clk => clk_0,
      nios2_clock_15_out_address_to_slave => nios2_clock_15_out_address_to_slave,
      nios2_clock_15_out_nativeaddress => nios2_clock_15_out_nativeaddress,
      nios2_clock_15_out_read => nios2_clock_15_out_read,
      nios2_clock_15_out_write => nios2_clock_15_out_write,
      nios2_clock_15_out_writedata => nios2_clock_15_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_cal_dac_code_pio, which is an e_ptf_instance
  the_cal_dac_code_pio : cal_dac_code_pio
    port map(
      out_port => internal_out_port_from_the_cal_dac_code_pio,
      readdata => cal_dac_code_pio_s1_readdata,
      address => cal_dac_code_pio_s1_address,
      chipselect => cal_dac_code_pio_s1_chipselect,
      clk => clk_0,
      reset_n => cal_dac_code_pio_s1_reset_n,
      write_n => cal_dac_code_pio_s1_write_n,
      writedata => cal_dac_code_pio_s1_writedata
    );


  --the_comparator_pio_s1, which is an e_instance
  the_comparator_pio_s1 : comparator_pio_s1_arbitrator
    port map(
      comparator_pio_s1_address => comparator_pio_s1_address,
      comparator_pio_s1_readdata_from_sa => comparator_pio_s1_readdata_from_sa,
      comparator_pio_s1_reset_n => comparator_pio_s1_reset_n,
      d1_comparator_pio_s1_end_xfer => d1_comparator_pio_s1_end_xfer,
      nios2_clock_11_out_granted_comparator_pio_s1 => nios2_clock_11_out_granted_comparator_pio_s1,
      nios2_clock_11_out_qualified_request_comparator_pio_s1 => nios2_clock_11_out_qualified_request_comparator_pio_s1,
      nios2_clock_11_out_read_data_valid_comparator_pio_s1 => nios2_clock_11_out_read_data_valid_comparator_pio_s1,
      nios2_clock_11_out_requests_comparator_pio_s1 => nios2_clock_11_out_requests_comparator_pio_s1,
      clk => internal_altpll_0_c0,
      comparator_pio_s1_readdata => comparator_pio_s1_readdata,
      nios2_clock_11_out_address_to_slave => nios2_clock_11_out_address_to_slave,
      nios2_clock_11_out_nativeaddress => nios2_clock_11_out_nativeaddress,
      nios2_clock_11_out_read => nios2_clock_11_out_read,
      nios2_clock_11_out_write => nios2_clock_11_out_write,
      reset_n => altpll_0_c0_reset_n
    );


  --the_comparator_pio, which is an e_ptf_instance
  the_comparator_pio : comparator_pio
    port map(
      readdata => comparator_pio_s1_readdata,
      address => comparator_pio_s1_address,
      clk => internal_altpll_0_c0,
      in_port => in_port_to_the_comparator_pio,
      reset_n => comparator_pio_s1_reset_n
    );


  --the_cpu_0_jtag_debug_module, which is an e_instance
  the_cpu_0_jtag_debug_module : cpu_0_jtag_debug_module_arbitrator
    port map(
      cpu_0_data_master_granted_cpu_0_jtag_debug_module => cpu_0_data_master_granted_cpu_0_jtag_debug_module,
      cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_data_master_requests_cpu_0_jtag_debug_module => cpu_0_data_master_requests_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_granted_cpu_0_jtag_debug_module => cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_requests_cpu_0_jtag_debug_module => cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
      cpu_0_jtag_debug_module_address => cpu_0_jtag_debug_module_address,
      cpu_0_jtag_debug_module_begintransfer => cpu_0_jtag_debug_module_begintransfer,
      cpu_0_jtag_debug_module_byteenable => cpu_0_jtag_debug_module_byteenable,
      cpu_0_jtag_debug_module_chipselect => cpu_0_jtag_debug_module_chipselect,
      cpu_0_jtag_debug_module_debugaccess => cpu_0_jtag_debug_module_debugaccess,
      cpu_0_jtag_debug_module_readdata_from_sa => cpu_0_jtag_debug_module_readdata_from_sa,
      cpu_0_jtag_debug_module_reset_n => cpu_0_jtag_debug_module_reset_n,
      cpu_0_jtag_debug_module_resetrequest_from_sa => cpu_0_jtag_debug_module_resetrequest_from_sa,
      cpu_0_jtag_debug_module_write => cpu_0_jtag_debug_module_write,
      cpu_0_jtag_debug_module_writedata => cpu_0_jtag_debug_module_writedata,
      d1_cpu_0_jtag_debug_module_end_xfer => d1_cpu_0_jtag_debug_module_end_xfer,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_debugaccess => cpu_0_data_master_debugaccess,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_latency_counter => cpu_0_instruction_master_latency_counter,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      cpu_0_jtag_debug_module_readdata => cpu_0_jtag_debug_module_readdata,
      cpu_0_jtag_debug_module_resetrequest => cpu_0_jtag_debug_module_resetrequest,
      reset_n => processor_clk_reset_n
    );


  --the_cpu_0_data_master, which is an e_instance
  the_cpu_0_data_master : cpu_0_data_master_arbitrator
    port map(
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_dbs_address => cpu_0_data_master_dbs_address,
      cpu_0_data_master_dbs_write_16 => cpu_0_data_master_dbs_write_16,
      cpu_0_data_master_irq => cpu_0_data_master_irq,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_readdata => cpu_0_data_master_readdata,
      cpu_0_data_master_readdatavalid => cpu_0_data_master_readdatavalid,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      clk => processor_clk,
      cpu_0_data_master_address => cpu_0_data_master_address,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_byteenable_nios2_clock_9_in => cpu_0_data_master_byteenable_nios2_clock_9_in,
      cpu_0_data_master_granted_cpu_0_jtag_debug_module => cpu_0_data_master_granted_cpu_0_jtag_debug_module,
      cpu_0_data_master_granted_nios2_clock_10_in => cpu_0_data_master_granted_nios2_clock_10_in,
      cpu_0_data_master_granted_nios2_clock_11_in => cpu_0_data_master_granted_nios2_clock_11_in,
      cpu_0_data_master_granted_nios2_clock_12_in => cpu_0_data_master_granted_nios2_clock_12_in,
      cpu_0_data_master_granted_nios2_clock_13_in => cpu_0_data_master_granted_nios2_clock_13_in,
      cpu_0_data_master_granted_nios2_clock_14_in => cpu_0_data_master_granted_nios2_clock_14_in,
      cpu_0_data_master_granted_nios2_clock_15_in => cpu_0_data_master_granted_nios2_clock_15_in,
      cpu_0_data_master_granted_nios2_clock_16_in => cpu_0_data_master_granted_nios2_clock_16_in,
      cpu_0_data_master_granted_nios2_clock_17_in => cpu_0_data_master_granted_nios2_clock_17_in,
      cpu_0_data_master_granted_nios2_clock_18_in => cpu_0_data_master_granted_nios2_clock_18_in,
      cpu_0_data_master_granted_nios2_clock_1_in => cpu_0_data_master_granted_nios2_clock_1_in,
      cpu_0_data_master_granted_nios2_clock_2_in => cpu_0_data_master_granted_nios2_clock_2_in,
      cpu_0_data_master_granted_nios2_clock_3_in => cpu_0_data_master_granted_nios2_clock_3_in,
      cpu_0_data_master_granted_nios2_clock_4_in => cpu_0_data_master_granted_nios2_clock_4_in,
      cpu_0_data_master_granted_nios2_clock_5_in => cpu_0_data_master_granted_nios2_clock_5_in,
      cpu_0_data_master_granted_nios2_clock_6_in => cpu_0_data_master_granted_nios2_clock_6_in,
      cpu_0_data_master_granted_nios2_clock_7_in => cpu_0_data_master_granted_nios2_clock_7_in,
      cpu_0_data_master_granted_nios2_clock_9_in => cpu_0_data_master_granted_nios2_clock_9_in,
      cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_data_master_qualified_request_nios2_clock_10_in => cpu_0_data_master_qualified_request_nios2_clock_10_in,
      cpu_0_data_master_qualified_request_nios2_clock_11_in => cpu_0_data_master_qualified_request_nios2_clock_11_in,
      cpu_0_data_master_qualified_request_nios2_clock_12_in => cpu_0_data_master_qualified_request_nios2_clock_12_in,
      cpu_0_data_master_qualified_request_nios2_clock_13_in => cpu_0_data_master_qualified_request_nios2_clock_13_in,
      cpu_0_data_master_qualified_request_nios2_clock_14_in => cpu_0_data_master_qualified_request_nios2_clock_14_in,
      cpu_0_data_master_qualified_request_nios2_clock_15_in => cpu_0_data_master_qualified_request_nios2_clock_15_in,
      cpu_0_data_master_qualified_request_nios2_clock_16_in => cpu_0_data_master_qualified_request_nios2_clock_16_in,
      cpu_0_data_master_qualified_request_nios2_clock_17_in => cpu_0_data_master_qualified_request_nios2_clock_17_in,
      cpu_0_data_master_qualified_request_nios2_clock_18_in => cpu_0_data_master_qualified_request_nios2_clock_18_in,
      cpu_0_data_master_qualified_request_nios2_clock_1_in => cpu_0_data_master_qualified_request_nios2_clock_1_in,
      cpu_0_data_master_qualified_request_nios2_clock_2_in => cpu_0_data_master_qualified_request_nios2_clock_2_in,
      cpu_0_data_master_qualified_request_nios2_clock_3_in => cpu_0_data_master_qualified_request_nios2_clock_3_in,
      cpu_0_data_master_qualified_request_nios2_clock_4_in => cpu_0_data_master_qualified_request_nios2_clock_4_in,
      cpu_0_data_master_qualified_request_nios2_clock_5_in => cpu_0_data_master_qualified_request_nios2_clock_5_in,
      cpu_0_data_master_qualified_request_nios2_clock_6_in => cpu_0_data_master_qualified_request_nios2_clock_6_in,
      cpu_0_data_master_qualified_request_nios2_clock_7_in => cpu_0_data_master_qualified_request_nios2_clock_7_in,
      cpu_0_data_master_qualified_request_nios2_clock_9_in => cpu_0_data_master_qualified_request_nios2_clock_9_in,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_data_master_read_data_valid_nios2_clock_10_in => cpu_0_data_master_read_data_valid_nios2_clock_10_in,
      cpu_0_data_master_read_data_valid_nios2_clock_11_in => cpu_0_data_master_read_data_valid_nios2_clock_11_in,
      cpu_0_data_master_read_data_valid_nios2_clock_12_in => cpu_0_data_master_read_data_valid_nios2_clock_12_in,
      cpu_0_data_master_read_data_valid_nios2_clock_13_in => cpu_0_data_master_read_data_valid_nios2_clock_13_in,
      cpu_0_data_master_read_data_valid_nios2_clock_14_in => cpu_0_data_master_read_data_valid_nios2_clock_14_in,
      cpu_0_data_master_read_data_valid_nios2_clock_15_in => cpu_0_data_master_read_data_valid_nios2_clock_15_in,
      cpu_0_data_master_read_data_valid_nios2_clock_16_in => cpu_0_data_master_read_data_valid_nios2_clock_16_in,
      cpu_0_data_master_read_data_valid_nios2_clock_17_in => cpu_0_data_master_read_data_valid_nios2_clock_17_in,
      cpu_0_data_master_read_data_valid_nios2_clock_18_in => cpu_0_data_master_read_data_valid_nios2_clock_18_in,
      cpu_0_data_master_read_data_valid_nios2_clock_1_in => cpu_0_data_master_read_data_valid_nios2_clock_1_in,
      cpu_0_data_master_read_data_valid_nios2_clock_2_in => cpu_0_data_master_read_data_valid_nios2_clock_2_in,
      cpu_0_data_master_read_data_valid_nios2_clock_3_in => cpu_0_data_master_read_data_valid_nios2_clock_3_in,
      cpu_0_data_master_read_data_valid_nios2_clock_4_in => cpu_0_data_master_read_data_valid_nios2_clock_4_in,
      cpu_0_data_master_read_data_valid_nios2_clock_5_in => cpu_0_data_master_read_data_valid_nios2_clock_5_in,
      cpu_0_data_master_read_data_valid_nios2_clock_6_in => cpu_0_data_master_read_data_valid_nios2_clock_6_in,
      cpu_0_data_master_read_data_valid_nios2_clock_7_in => cpu_0_data_master_read_data_valid_nios2_clock_7_in,
      cpu_0_data_master_read_data_valid_nios2_clock_9_in => cpu_0_data_master_read_data_valid_nios2_clock_9_in,
      cpu_0_data_master_requests_cpu_0_jtag_debug_module => cpu_0_data_master_requests_cpu_0_jtag_debug_module,
      cpu_0_data_master_requests_nios2_clock_10_in => cpu_0_data_master_requests_nios2_clock_10_in,
      cpu_0_data_master_requests_nios2_clock_11_in => cpu_0_data_master_requests_nios2_clock_11_in,
      cpu_0_data_master_requests_nios2_clock_12_in => cpu_0_data_master_requests_nios2_clock_12_in,
      cpu_0_data_master_requests_nios2_clock_13_in => cpu_0_data_master_requests_nios2_clock_13_in,
      cpu_0_data_master_requests_nios2_clock_14_in => cpu_0_data_master_requests_nios2_clock_14_in,
      cpu_0_data_master_requests_nios2_clock_15_in => cpu_0_data_master_requests_nios2_clock_15_in,
      cpu_0_data_master_requests_nios2_clock_16_in => cpu_0_data_master_requests_nios2_clock_16_in,
      cpu_0_data_master_requests_nios2_clock_17_in => cpu_0_data_master_requests_nios2_clock_17_in,
      cpu_0_data_master_requests_nios2_clock_18_in => cpu_0_data_master_requests_nios2_clock_18_in,
      cpu_0_data_master_requests_nios2_clock_1_in => cpu_0_data_master_requests_nios2_clock_1_in,
      cpu_0_data_master_requests_nios2_clock_2_in => cpu_0_data_master_requests_nios2_clock_2_in,
      cpu_0_data_master_requests_nios2_clock_3_in => cpu_0_data_master_requests_nios2_clock_3_in,
      cpu_0_data_master_requests_nios2_clock_4_in => cpu_0_data_master_requests_nios2_clock_4_in,
      cpu_0_data_master_requests_nios2_clock_5_in => cpu_0_data_master_requests_nios2_clock_5_in,
      cpu_0_data_master_requests_nios2_clock_6_in => cpu_0_data_master_requests_nios2_clock_6_in,
      cpu_0_data_master_requests_nios2_clock_7_in => cpu_0_data_master_requests_nios2_clock_7_in,
      cpu_0_data_master_requests_nios2_clock_9_in => cpu_0_data_master_requests_nios2_clock_9_in,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      cpu_0_jtag_debug_module_readdata_from_sa => cpu_0_jtag_debug_module_readdata_from_sa,
      d1_cpu_0_jtag_debug_module_end_xfer => d1_cpu_0_jtag_debug_module_end_xfer,
      d1_nios2_clock_10_in_end_xfer => d1_nios2_clock_10_in_end_xfer,
      d1_nios2_clock_11_in_end_xfer => d1_nios2_clock_11_in_end_xfer,
      d1_nios2_clock_12_in_end_xfer => d1_nios2_clock_12_in_end_xfer,
      d1_nios2_clock_13_in_end_xfer => d1_nios2_clock_13_in_end_xfer,
      d1_nios2_clock_14_in_end_xfer => d1_nios2_clock_14_in_end_xfer,
      d1_nios2_clock_15_in_end_xfer => d1_nios2_clock_15_in_end_xfer,
      d1_nios2_clock_16_in_end_xfer => d1_nios2_clock_16_in_end_xfer,
      d1_nios2_clock_17_in_end_xfer => d1_nios2_clock_17_in_end_xfer,
      d1_nios2_clock_18_in_end_xfer => d1_nios2_clock_18_in_end_xfer,
      d1_nios2_clock_1_in_end_xfer => d1_nios2_clock_1_in_end_xfer,
      d1_nios2_clock_2_in_end_xfer => d1_nios2_clock_2_in_end_xfer,
      d1_nios2_clock_3_in_end_xfer => d1_nios2_clock_3_in_end_xfer,
      d1_nios2_clock_4_in_end_xfer => d1_nios2_clock_4_in_end_xfer,
      d1_nios2_clock_5_in_end_xfer => d1_nios2_clock_5_in_end_xfer,
      d1_nios2_clock_6_in_end_xfer => d1_nios2_clock_6_in_end_xfer,
      d1_nios2_clock_7_in_end_xfer => d1_nios2_clock_7_in_end_xfer,
      d1_nios2_clock_9_in_end_xfer => d1_nios2_clock_9_in_end_xfer,
      jtag_uart_0_avalon_jtag_slave_irq_from_sa => jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      nios2_clock_10_in_readdata_from_sa => nios2_clock_10_in_readdata_from_sa,
      nios2_clock_10_in_waitrequest_from_sa => nios2_clock_10_in_waitrequest_from_sa,
      nios2_clock_11_in_readdata_from_sa => nios2_clock_11_in_readdata_from_sa,
      nios2_clock_11_in_waitrequest_from_sa => nios2_clock_11_in_waitrequest_from_sa,
      nios2_clock_12_in_readdata_from_sa => nios2_clock_12_in_readdata_from_sa,
      nios2_clock_12_in_waitrequest_from_sa => nios2_clock_12_in_waitrequest_from_sa,
      nios2_clock_13_in_readdata_from_sa => nios2_clock_13_in_readdata_from_sa,
      nios2_clock_13_in_waitrequest_from_sa => nios2_clock_13_in_waitrequest_from_sa,
      nios2_clock_14_in_readdata_from_sa => nios2_clock_14_in_readdata_from_sa,
      nios2_clock_14_in_waitrequest_from_sa => nios2_clock_14_in_waitrequest_from_sa,
      nios2_clock_15_in_readdata_from_sa => nios2_clock_15_in_readdata_from_sa,
      nios2_clock_15_in_waitrequest_from_sa => nios2_clock_15_in_waitrequest_from_sa,
      nios2_clock_16_in_readdata_from_sa => nios2_clock_16_in_readdata_from_sa,
      nios2_clock_16_in_waitrequest_from_sa => nios2_clock_16_in_waitrequest_from_sa,
      nios2_clock_17_in_readdata_from_sa => nios2_clock_17_in_readdata_from_sa,
      nios2_clock_17_in_waitrequest_from_sa => nios2_clock_17_in_waitrequest_from_sa,
      nios2_clock_18_in_readdata_from_sa => nios2_clock_18_in_readdata_from_sa,
      nios2_clock_18_in_waitrequest_from_sa => nios2_clock_18_in_waitrequest_from_sa,
      nios2_clock_1_in_readdata_from_sa => nios2_clock_1_in_readdata_from_sa,
      nios2_clock_1_in_waitrequest_from_sa => nios2_clock_1_in_waitrequest_from_sa,
      nios2_clock_2_in_readdata_from_sa => nios2_clock_2_in_readdata_from_sa,
      nios2_clock_2_in_waitrequest_from_sa => nios2_clock_2_in_waitrequest_from_sa,
      nios2_clock_3_in_readdata_from_sa => nios2_clock_3_in_readdata_from_sa,
      nios2_clock_3_in_waitrequest_from_sa => nios2_clock_3_in_waitrequest_from_sa,
      nios2_clock_4_in_readdata_from_sa => nios2_clock_4_in_readdata_from_sa,
      nios2_clock_4_in_waitrequest_from_sa => nios2_clock_4_in_waitrequest_from_sa,
      nios2_clock_5_in_readdata_from_sa => nios2_clock_5_in_readdata_from_sa,
      nios2_clock_5_in_waitrequest_from_sa => nios2_clock_5_in_waitrequest_from_sa,
      nios2_clock_6_in_readdata_from_sa => nios2_clock_6_in_readdata_from_sa,
      nios2_clock_6_in_waitrequest_from_sa => nios2_clock_6_in_waitrequest_from_sa,
      nios2_clock_7_in_readdata_from_sa => nios2_clock_7_in_readdata_from_sa,
      nios2_clock_7_in_waitrequest_from_sa => nios2_clock_7_in_waitrequest_from_sa,
      nios2_clock_9_in_readdata_from_sa => nios2_clock_9_in_readdata_from_sa,
      nios2_clock_9_in_waitrequest_from_sa => nios2_clock_9_in_waitrequest_from_sa,
      processor_clk => processor_clk,
      processor_clk_reset_n => processor_clk_reset_n,
      reset_n => processor_clk_reset_n,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa
    );


  --the_cpu_0_instruction_master, which is an e_instance
  the_cpu_0_instruction_master : cpu_0_instruction_master_arbitrator
    port map(
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_dbs_address => cpu_0_instruction_master_dbs_address,
      cpu_0_instruction_master_latency_counter => cpu_0_instruction_master_latency_counter,
      cpu_0_instruction_master_readdata => cpu_0_instruction_master_readdata,
      cpu_0_instruction_master_readdatavalid => cpu_0_instruction_master_readdatavalid,
      cpu_0_instruction_master_waitrequest => cpu_0_instruction_master_waitrequest,
      clk => processor_clk,
      cpu_0_instruction_master_address => cpu_0_instruction_master_address,
      cpu_0_instruction_master_granted_cpu_0_jtag_debug_module => cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_granted_nios2_clock_0_in => cpu_0_instruction_master_granted_nios2_clock_0_in,
      cpu_0_instruction_master_granted_nios2_clock_8_in => cpu_0_instruction_master_granted_nios2_clock_8_in,
      cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_qualified_request_nios2_clock_0_in => cpu_0_instruction_master_qualified_request_nios2_clock_0_in,
      cpu_0_instruction_master_qualified_request_nios2_clock_8_in => cpu_0_instruction_master_qualified_request_nios2_clock_8_in,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_read_data_valid_nios2_clock_0_in => cpu_0_instruction_master_read_data_valid_nios2_clock_0_in,
      cpu_0_instruction_master_read_data_valid_nios2_clock_8_in => cpu_0_instruction_master_read_data_valid_nios2_clock_8_in,
      cpu_0_instruction_master_requests_cpu_0_jtag_debug_module => cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_requests_nios2_clock_0_in => cpu_0_instruction_master_requests_nios2_clock_0_in,
      cpu_0_instruction_master_requests_nios2_clock_8_in => cpu_0_instruction_master_requests_nios2_clock_8_in,
      cpu_0_jtag_debug_module_readdata_from_sa => cpu_0_jtag_debug_module_readdata_from_sa,
      d1_cpu_0_jtag_debug_module_end_xfer => d1_cpu_0_jtag_debug_module_end_xfer,
      d1_nios2_clock_0_in_end_xfer => d1_nios2_clock_0_in_end_xfer,
      d1_nios2_clock_8_in_end_xfer => d1_nios2_clock_8_in_end_xfer,
      nios2_clock_0_in_readdata_from_sa => nios2_clock_0_in_readdata_from_sa,
      nios2_clock_0_in_waitrequest_from_sa => nios2_clock_0_in_waitrequest_from_sa,
      nios2_clock_8_in_readdata_from_sa => nios2_clock_8_in_readdata_from_sa,
      nios2_clock_8_in_waitrequest_from_sa => nios2_clock_8_in_waitrequest_from_sa,
      reset_n => processor_clk_reset_n
    );


  --the_cpu_0, which is an e_ptf_instance
  the_cpu_0 : cpu_0
    port map(
      d_address => cpu_0_data_master_address,
      d_byteenable => cpu_0_data_master_byteenable,
      d_read => cpu_0_data_master_read,
      d_write => cpu_0_data_master_write,
      d_writedata => cpu_0_data_master_writedata,
      i_address => cpu_0_instruction_master_address,
      i_read => cpu_0_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => cpu_0_data_master_debugaccess,
      jtag_debug_module_readdata => cpu_0_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => cpu_0_jtag_debug_module_resetrequest,
      clk => processor_clk,
      d_irq => cpu_0_data_master_irq,
      d_readdata => cpu_0_data_master_readdata,
      d_readdatavalid => cpu_0_data_master_readdatavalid,
      d_waitrequest => cpu_0_data_master_waitrequest,
      i_readdata => cpu_0_instruction_master_readdata,
      i_readdatavalid => cpu_0_instruction_master_readdatavalid,
      i_waitrequest => cpu_0_instruction_master_waitrequest,
      jtag_debug_module_address => cpu_0_jtag_debug_module_address,
      jtag_debug_module_begintransfer => cpu_0_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => cpu_0_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => cpu_0_jtag_debug_module_debugaccess,
      jtag_debug_module_select => cpu_0_jtag_debug_module_chipselect,
      jtag_debug_module_write => cpu_0_jtag_debug_module_write,
      jtag_debug_module_writedata => cpu_0_jtag_debug_module_writedata,
      reset_n => cpu_0_jtag_debug_module_reset_n
    );


  --the_gen_code_strobe_s1, which is an e_instance
  the_gen_code_strobe_s1 : gen_code_strobe_s1_arbitrator
    port map(
      d1_gen_code_strobe_s1_end_xfer => d1_gen_code_strobe_s1_end_xfer,
      gen_code_strobe_s1_address => gen_code_strobe_s1_address,
      gen_code_strobe_s1_chipselect => gen_code_strobe_s1_chipselect,
      gen_code_strobe_s1_readdata_from_sa => gen_code_strobe_s1_readdata_from_sa,
      gen_code_strobe_s1_reset_n => gen_code_strobe_s1_reset_n,
      gen_code_strobe_s1_write_n => gen_code_strobe_s1_write_n,
      gen_code_strobe_s1_writedata => gen_code_strobe_s1_writedata,
      nios2_clock_13_out_granted_gen_code_strobe_s1 => nios2_clock_13_out_granted_gen_code_strobe_s1,
      nios2_clock_13_out_qualified_request_gen_code_strobe_s1 => nios2_clock_13_out_qualified_request_gen_code_strobe_s1,
      nios2_clock_13_out_read_data_valid_gen_code_strobe_s1 => nios2_clock_13_out_read_data_valid_gen_code_strobe_s1,
      nios2_clock_13_out_requests_gen_code_strobe_s1 => nios2_clock_13_out_requests_gen_code_strobe_s1,
      clk => clk_0,
      gen_code_strobe_s1_readdata => gen_code_strobe_s1_readdata,
      nios2_clock_13_out_address_to_slave => nios2_clock_13_out_address_to_slave,
      nios2_clock_13_out_nativeaddress => nios2_clock_13_out_nativeaddress,
      nios2_clock_13_out_read => nios2_clock_13_out_read,
      nios2_clock_13_out_write => nios2_clock_13_out_write,
      nios2_clock_13_out_writedata => nios2_clock_13_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_gen_code_strobe, which is an e_ptf_instance
  the_gen_code_strobe : gen_code_strobe
    port map(
      out_port => internal_out_port_from_the_gen_code_strobe,
      readdata => gen_code_strobe_s1_readdata,
      address => gen_code_strobe_s1_address,
      chipselect => gen_code_strobe_s1_chipselect,
      clk => clk_0,
      reset_n => gen_code_strobe_s1_reset_n,
      write_n => gen_code_strobe_s1_write_n,
      writedata => gen_code_strobe_s1_writedata
    );


  --the_gen_code_value_pio_0_s1, which is an e_instance
  the_gen_code_value_pio_0_s1 : gen_code_value_pio_0_s1_arbitrator
    port map(
      d1_gen_code_value_pio_0_s1_end_xfer => d1_gen_code_value_pio_0_s1_end_xfer,
      gen_code_value_pio_0_s1_address => gen_code_value_pio_0_s1_address,
      gen_code_value_pio_0_s1_chipselect => gen_code_value_pio_0_s1_chipselect,
      gen_code_value_pio_0_s1_readdata_from_sa => gen_code_value_pio_0_s1_readdata_from_sa,
      gen_code_value_pio_0_s1_reset_n => gen_code_value_pio_0_s1_reset_n,
      gen_code_value_pio_0_s1_write_n => gen_code_value_pio_0_s1_write_n,
      gen_code_value_pio_0_s1_writedata => gen_code_value_pio_0_s1_writedata,
      nios2_clock_6_out_granted_gen_code_value_pio_0_s1 => nios2_clock_6_out_granted_gen_code_value_pio_0_s1,
      nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 => nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1,
      nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1 => nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1,
      nios2_clock_6_out_requests_gen_code_value_pio_0_s1 => nios2_clock_6_out_requests_gen_code_value_pio_0_s1,
      clk => internal_altpll_0_c0,
      gen_code_value_pio_0_s1_readdata => gen_code_value_pio_0_s1_readdata,
      nios2_clock_6_out_address_to_slave => nios2_clock_6_out_address_to_slave,
      nios2_clock_6_out_nativeaddress => nios2_clock_6_out_nativeaddress,
      nios2_clock_6_out_read => nios2_clock_6_out_read,
      nios2_clock_6_out_write => nios2_clock_6_out_write,
      nios2_clock_6_out_writedata => nios2_clock_6_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_gen_code_value_pio_0, which is an e_ptf_instance
  the_gen_code_value_pio_0 : gen_code_value_pio_0
    port map(
      out_port => internal_out_port_from_the_gen_code_value_pio_0,
      readdata => gen_code_value_pio_0_s1_readdata,
      address => gen_code_value_pio_0_s1_address,
      chipselect => gen_code_value_pio_0_s1_chipselect,
      clk => internal_altpll_0_c0,
      reset_n => gen_code_value_pio_0_s1_reset_n,
      write_n => gen_code_value_pio_0_s1_write_n,
      writedata => gen_code_value_pio_0_s1_writedata
    );


  --the_gen_code_value_pio_1_s1, which is an e_instance
  the_gen_code_value_pio_1_s1 : gen_code_value_pio_1_s1_arbitrator
    port map(
      d1_gen_code_value_pio_1_s1_end_xfer => d1_gen_code_value_pio_1_s1_end_xfer,
      gen_code_value_pio_1_s1_address => gen_code_value_pio_1_s1_address,
      gen_code_value_pio_1_s1_chipselect => gen_code_value_pio_1_s1_chipselect,
      gen_code_value_pio_1_s1_readdata_from_sa => gen_code_value_pio_1_s1_readdata_from_sa,
      gen_code_value_pio_1_s1_reset_n => gen_code_value_pio_1_s1_reset_n,
      gen_code_value_pio_1_s1_write_n => gen_code_value_pio_1_s1_write_n,
      gen_code_value_pio_1_s1_writedata => gen_code_value_pio_1_s1_writedata,
      nios2_clock_7_out_granted_gen_code_value_pio_1_s1 => nios2_clock_7_out_granted_gen_code_value_pio_1_s1,
      nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 => nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1,
      nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1 => nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1,
      nios2_clock_7_out_requests_gen_code_value_pio_1_s1 => nios2_clock_7_out_requests_gen_code_value_pio_1_s1,
      clk => internal_altpll_0_c0,
      gen_code_value_pio_1_s1_readdata => gen_code_value_pio_1_s1_readdata,
      nios2_clock_7_out_address_to_slave => nios2_clock_7_out_address_to_slave,
      nios2_clock_7_out_nativeaddress => nios2_clock_7_out_nativeaddress,
      nios2_clock_7_out_read => nios2_clock_7_out_read,
      nios2_clock_7_out_write => nios2_clock_7_out_write,
      nios2_clock_7_out_writedata => nios2_clock_7_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_gen_code_value_pio_1, which is an e_ptf_instance
  the_gen_code_value_pio_1 : gen_code_value_pio_1
    port map(
      out_port => internal_out_port_from_the_gen_code_value_pio_1,
      readdata => gen_code_value_pio_1_s1_readdata,
      address => gen_code_value_pio_1_s1_address,
      chipselect => gen_code_value_pio_1_s1_chipselect,
      clk => internal_altpll_0_c0,
      reset_n => gen_code_value_pio_1_s1_reset_n,
      write_n => gen_code_value_pio_1_s1_write_n,
      writedata => gen_code_value_pio_1_s1_writedata
    );


  --the_jtag_uart_0_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_0_avalon_jtag_slave : jtag_uart_0_avalon_jtag_slave_arbitrator
    port map(
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer => d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
      jtag_uart_0_avalon_jtag_slave_address => jtag_uart_0_avalon_jtag_slave_address,
      jtag_uart_0_avalon_jtag_slave_chipselect => jtag_uart_0_avalon_jtag_slave_chipselect,
      jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_0_avalon_jtag_slave_irq_from_sa => jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      jtag_uart_0_avalon_jtag_slave_read_n => jtag_uart_0_avalon_jtag_slave_read_n,
      jtag_uart_0_avalon_jtag_slave_readdata_from_sa => jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_0_avalon_jtag_slave_reset_n => jtag_uart_0_avalon_jtag_slave_reset_n,
      jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_0_avalon_jtag_slave_write_n => jtag_uart_0_avalon_jtag_slave_write_n,
      jtag_uart_0_avalon_jtag_slave_writedata => jtag_uart_0_avalon_jtag_slave_writedata,
      nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave,
      nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave,
      nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave,
      nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave,
      clk => internal_altpll_0_c0,
      jtag_uart_0_avalon_jtag_slave_dataavailable => jtag_uart_0_avalon_jtag_slave_dataavailable,
      jtag_uart_0_avalon_jtag_slave_irq => jtag_uart_0_avalon_jtag_slave_irq,
      jtag_uart_0_avalon_jtag_slave_readdata => jtag_uart_0_avalon_jtag_slave_readdata,
      jtag_uart_0_avalon_jtag_slave_readyfordata => jtag_uart_0_avalon_jtag_slave_readyfordata,
      jtag_uart_0_avalon_jtag_slave_waitrequest => jtag_uart_0_avalon_jtag_slave_waitrequest,
      nios2_clock_2_out_address_to_slave => nios2_clock_2_out_address_to_slave,
      nios2_clock_2_out_nativeaddress => nios2_clock_2_out_nativeaddress,
      nios2_clock_2_out_read => nios2_clock_2_out_read,
      nios2_clock_2_out_write => nios2_clock_2_out_write,
      nios2_clock_2_out_writedata => nios2_clock_2_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_jtag_uart_0, which is an e_ptf_instance
  the_jtag_uart_0 : jtag_uart_0
    port map(
      av_irq => jtag_uart_0_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_0_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_0_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_0_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_0_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_0_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_0_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_0_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_0_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_0_avalon_jtag_slave_writedata,
      clk => internal_altpll_0_c0,
      rst_n => jtag_uart_0_avalon_jtag_slave_reset_n
    );


  --the_latch_pio_s1, which is an e_instance
  the_latch_pio_s1 : latch_pio_s1_arbitrator
    port map(
      d1_latch_pio_s1_end_xfer => d1_latch_pio_s1_end_xfer,
      latch_pio_s1_address => latch_pio_s1_address,
      latch_pio_s1_chipselect => latch_pio_s1_chipselect,
      latch_pio_s1_readdata_from_sa => latch_pio_s1_readdata_from_sa,
      latch_pio_s1_reset_n => latch_pio_s1_reset_n,
      latch_pio_s1_write_n => latch_pio_s1_write_n,
      latch_pio_s1_writedata => latch_pio_s1_writedata,
      nios2_clock_18_out_granted_latch_pio_s1 => nios2_clock_18_out_granted_latch_pio_s1,
      nios2_clock_18_out_qualified_request_latch_pio_s1 => nios2_clock_18_out_qualified_request_latch_pio_s1,
      nios2_clock_18_out_read_data_valid_latch_pio_s1 => nios2_clock_18_out_read_data_valid_latch_pio_s1,
      nios2_clock_18_out_requests_latch_pio_s1 => nios2_clock_18_out_requests_latch_pio_s1,
      clk => clk_0,
      latch_pio_s1_readdata => latch_pio_s1_readdata,
      nios2_clock_18_out_address_to_slave => nios2_clock_18_out_address_to_slave,
      nios2_clock_18_out_nativeaddress => nios2_clock_18_out_nativeaddress,
      nios2_clock_18_out_read => nios2_clock_18_out_read,
      nios2_clock_18_out_write => nios2_clock_18_out_write,
      nios2_clock_18_out_writedata => nios2_clock_18_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_latch_pio, which is an e_ptf_instance
  the_latch_pio : latch_pio
    port map(
      out_port => internal_out_port_from_the_latch_pio,
      readdata => latch_pio_s1_readdata,
      address => latch_pio_s1_address,
      chipselect => latch_pio_s1_chipselect,
      clk => clk_0,
      reset_n => latch_pio_s1_reset_n,
      write_n => latch_pio_s1_write_n,
      writedata => latch_pio_s1_writedata
    );


  --the_led_pio_s1, which is an e_instance
  the_led_pio_s1 : led_pio_s1_arbitrator
    port map(
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      led_pio_s1_address => led_pio_s1_address,
      led_pio_s1_chipselect => led_pio_s1_chipselect,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      led_pio_s1_reset_n => led_pio_s1_reset_n,
      led_pio_s1_write_n => led_pio_s1_write_n,
      led_pio_s1_writedata => led_pio_s1_writedata,
      nios2_clock_12_out_granted_led_pio_s1 => nios2_clock_12_out_granted_led_pio_s1,
      nios2_clock_12_out_qualified_request_led_pio_s1 => nios2_clock_12_out_qualified_request_led_pio_s1,
      nios2_clock_12_out_read_data_valid_led_pio_s1 => nios2_clock_12_out_read_data_valid_led_pio_s1,
      nios2_clock_12_out_requests_led_pio_s1 => nios2_clock_12_out_requests_led_pio_s1,
      clk => clk_0,
      led_pio_s1_readdata => led_pio_s1_readdata,
      nios2_clock_12_out_address_to_slave => nios2_clock_12_out_address_to_slave,
      nios2_clock_12_out_nativeaddress => nios2_clock_12_out_nativeaddress,
      nios2_clock_12_out_read => nios2_clock_12_out_read,
      nios2_clock_12_out_write => nios2_clock_12_out_write,
      nios2_clock_12_out_writedata => nios2_clock_12_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_led_pio, which is an e_ptf_instance
  the_led_pio : led_pio
    port map(
      out_port => internal_out_port_from_the_led_pio,
      readdata => led_pio_s1_readdata,
      address => led_pio_s1_address,
      chipselect => led_pio_s1_chipselect,
      clk => clk_0,
      reset_n => led_pio_s1_reset_n,
      write_n => led_pio_s1_write_n,
      writedata => led_pio_s1_writedata
    );


  --the_mode_select_s1, which is an e_instance
  the_mode_select_s1 : mode_select_s1_arbitrator
    port map(
      d1_mode_select_s1_end_xfer => d1_mode_select_s1_end_xfer,
      mode_select_s1_address => mode_select_s1_address,
      mode_select_s1_chipselect => mode_select_s1_chipselect,
      mode_select_s1_readdata_from_sa => mode_select_s1_readdata_from_sa,
      mode_select_s1_reset_n => mode_select_s1_reset_n,
      mode_select_s1_write_n => mode_select_s1_write_n,
      mode_select_s1_writedata => mode_select_s1_writedata,
      nios2_clock_10_out_granted_mode_select_s1 => nios2_clock_10_out_granted_mode_select_s1,
      nios2_clock_10_out_qualified_request_mode_select_s1 => nios2_clock_10_out_qualified_request_mode_select_s1,
      nios2_clock_10_out_read_data_valid_mode_select_s1 => nios2_clock_10_out_read_data_valid_mode_select_s1,
      nios2_clock_10_out_requests_mode_select_s1 => nios2_clock_10_out_requests_mode_select_s1,
      clk => internal_altpll_0_c0,
      mode_select_s1_readdata => mode_select_s1_readdata,
      nios2_clock_10_out_address_to_slave => nios2_clock_10_out_address_to_slave,
      nios2_clock_10_out_nativeaddress => nios2_clock_10_out_nativeaddress,
      nios2_clock_10_out_read => nios2_clock_10_out_read,
      nios2_clock_10_out_write => nios2_clock_10_out_write,
      nios2_clock_10_out_writedata => nios2_clock_10_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_mode_select, which is an e_ptf_instance
  the_mode_select : mode_select
    port map(
      readdata => mode_select_s1_readdata,
      address => mode_select_s1_address,
      chipselect => mode_select_s1_chipselect,
      clk => internal_altpll_0_c0,
      in_port => in_port_to_the_mode_select,
      reset_n => mode_select_s1_reset_n,
      write_n => mode_select_s1_write_n,
      writedata => mode_select_s1_writedata
    );


  --the_nios2_clock_0_in, which is an e_instance
  the_nios2_clock_0_in : nios2_clock_0_in_arbitrator
    port map(
      cpu_0_instruction_master_granted_nios2_clock_0_in => cpu_0_instruction_master_granted_nios2_clock_0_in,
      cpu_0_instruction_master_qualified_request_nios2_clock_0_in => cpu_0_instruction_master_qualified_request_nios2_clock_0_in,
      cpu_0_instruction_master_read_data_valid_nios2_clock_0_in => cpu_0_instruction_master_read_data_valid_nios2_clock_0_in,
      cpu_0_instruction_master_requests_nios2_clock_0_in => cpu_0_instruction_master_requests_nios2_clock_0_in,
      d1_nios2_clock_0_in_end_xfer => d1_nios2_clock_0_in_end_xfer,
      nios2_clock_0_in_address => nios2_clock_0_in_address,
      nios2_clock_0_in_byteenable => nios2_clock_0_in_byteenable,
      nios2_clock_0_in_endofpacket_from_sa => nios2_clock_0_in_endofpacket_from_sa,
      nios2_clock_0_in_nativeaddress => nios2_clock_0_in_nativeaddress,
      nios2_clock_0_in_read => nios2_clock_0_in_read,
      nios2_clock_0_in_readdata_from_sa => nios2_clock_0_in_readdata_from_sa,
      nios2_clock_0_in_reset_n => nios2_clock_0_in_reset_n,
      nios2_clock_0_in_waitrequest_from_sa => nios2_clock_0_in_waitrequest_from_sa,
      nios2_clock_0_in_write => nios2_clock_0_in_write,
      clk => processor_clk,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_latency_counter => cpu_0_instruction_master_latency_counter,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      nios2_clock_0_in_endofpacket => nios2_clock_0_in_endofpacket,
      nios2_clock_0_in_readdata => nios2_clock_0_in_readdata,
      nios2_clock_0_in_waitrequest => nios2_clock_0_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_0_out, which is an e_instance
  the_nios2_clock_0_out : nios2_clock_0_out_arbitrator
    port map(
      nios2_clock_0_out_address_to_slave => nios2_clock_0_out_address_to_slave,
      nios2_clock_0_out_readdata => nios2_clock_0_out_readdata,
      nios2_clock_0_out_reset_n => nios2_clock_0_out_reset_n,
      nios2_clock_0_out_waitrequest => nios2_clock_0_out_waitrequest,
      clk => internal_altpll_0_c0,
      d1_onchip_mem_s1_end_xfer => d1_onchip_mem_s1_end_xfer,
      nios2_clock_0_out_address => nios2_clock_0_out_address,
      nios2_clock_0_out_byteenable => nios2_clock_0_out_byteenable,
      nios2_clock_0_out_granted_onchip_mem_s1 => nios2_clock_0_out_granted_onchip_mem_s1,
      nios2_clock_0_out_qualified_request_onchip_mem_s1 => nios2_clock_0_out_qualified_request_onchip_mem_s1,
      nios2_clock_0_out_read => nios2_clock_0_out_read,
      nios2_clock_0_out_read_data_valid_onchip_mem_s1 => nios2_clock_0_out_read_data_valid_onchip_mem_s1,
      nios2_clock_0_out_requests_onchip_mem_s1 => nios2_clock_0_out_requests_onchip_mem_s1,
      nios2_clock_0_out_write => nios2_clock_0_out_write,
      nios2_clock_0_out_writedata => nios2_clock_0_out_writedata,
      onchip_mem_s1_readdata_from_sa => onchip_mem_s1_readdata_from_sa,
      reset_n => altpll_0_c0_reset_n
    );


  --the_nios2_clock_0, which is an e_ptf_instance
  the_nios2_clock_0 : nios2_clock_0
    port map(
      master_address => nios2_clock_0_out_address,
      master_byteenable => nios2_clock_0_out_byteenable,
      master_nativeaddress => nios2_clock_0_out_nativeaddress,
      master_read => nios2_clock_0_out_read,
      master_write => nios2_clock_0_out_write,
      master_writedata => nios2_clock_0_out_writedata,
      slave_endofpacket => nios2_clock_0_in_endofpacket,
      slave_readdata => nios2_clock_0_in_readdata,
      slave_waitrequest => nios2_clock_0_in_waitrequest,
      master_clk => internal_altpll_0_c0,
      master_endofpacket => nios2_clock_0_out_endofpacket,
      master_readdata => nios2_clock_0_out_readdata,
      master_reset_n => nios2_clock_0_out_reset_n,
      master_waitrequest => nios2_clock_0_out_waitrequest,
      slave_address => nios2_clock_0_in_address,
      slave_byteenable => nios2_clock_0_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_0_in_nativeaddress,
      slave_read => nios2_clock_0_in_read,
      slave_reset_n => nios2_clock_0_in_reset_n,
      slave_write => nios2_clock_0_in_write,
      slave_writedata => nios2_clock_0_in_writedata
    );


  --the_nios2_clock_1_in, which is an e_instance
  the_nios2_clock_1_in : nios2_clock_1_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_1_in => cpu_0_data_master_granted_nios2_clock_1_in,
      cpu_0_data_master_qualified_request_nios2_clock_1_in => cpu_0_data_master_qualified_request_nios2_clock_1_in,
      cpu_0_data_master_read_data_valid_nios2_clock_1_in => cpu_0_data_master_read_data_valid_nios2_clock_1_in,
      cpu_0_data_master_requests_nios2_clock_1_in => cpu_0_data_master_requests_nios2_clock_1_in,
      d1_nios2_clock_1_in_end_xfer => d1_nios2_clock_1_in_end_xfer,
      nios2_clock_1_in_address => nios2_clock_1_in_address,
      nios2_clock_1_in_byteenable => nios2_clock_1_in_byteenable,
      nios2_clock_1_in_endofpacket_from_sa => nios2_clock_1_in_endofpacket_from_sa,
      nios2_clock_1_in_nativeaddress => nios2_clock_1_in_nativeaddress,
      nios2_clock_1_in_read => nios2_clock_1_in_read,
      nios2_clock_1_in_readdata_from_sa => nios2_clock_1_in_readdata_from_sa,
      nios2_clock_1_in_reset_n => nios2_clock_1_in_reset_n,
      nios2_clock_1_in_waitrequest_from_sa => nios2_clock_1_in_waitrequest_from_sa,
      nios2_clock_1_in_write => nios2_clock_1_in_write,
      nios2_clock_1_in_writedata => nios2_clock_1_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_1_in_endofpacket => nios2_clock_1_in_endofpacket,
      nios2_clock_1_in_readdata => nios2_clock_1_in_readdata,
      nios2_clock_1_in_waitrequest => nios2_clock_1_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_1_out, which is an e_instance
  the_nios2_clock_1_out : nios2_clock_1_out_arbitrator
    port map(
      nios2_clock_1_out_address_to_slave => nios2_clock_1_out_address_to_slave,
      nios2_clock_1_out_readdata => nios2_clock_1_out_readdata,
      nios2_clock_1_out_reset_n => nios2_clock_1_out_reset_n,
      nios2_clock_1_out_waitrequest => nios2_clock_1_out_waitrequest,
      clk => internal_altpll_0_c0,
      d1_onchip_mem_s1_end_xfer => d1_onchip_mem_s1_end_xfer,
      nios2_clock_1_out_address => nios2_clock_1_out_address,
      nios2_clock_1_out_byteenable => nios2_clock_1_out_byteenable,
      nios2_clock_1_out_granted_onchip_mem_s1 => nios2_clock_1_out_granted_onchip_mem_s1,
      nios2_clock_1_out_qualified_request_onchip_mem_s1 => nios2_clock_1_out_qualified_request_onchip_mem_s1,
      nios2_clock_1_out_read => nios2_clock_1_out_read,
      nios2_clock_1_out_read_data_valid_onchip_mem_s1 => nios2_clock_1_out_read_data_valid_onchip_mem_s1,
      nios2_clock_1_out_requests_onchip_mem_s1 => nios2_clock_1_out_requests_onchip_mem_s1,
      nios2_clock_1_out_write => nios2_clock_1_out_write,
      nios2_clock_1_out_writedata => nios2_clock_1_out_writedata,
      onchip_mem_s1_readdata_from_sa => onchip_mem_s1_readdata_from_sa,
      reset_n => altpll_0_c0_reset_n
    );


  --the_nios2_clock_1, which is an e_ptf_instance
  the_nios2_clock_1 : nios2_clock_1
    port map(
      master_address => nios2_clock_1_out_address,
      master_byteenable => nios2_clock_1_out_byteenable,
      master_nativeaddress => nios2_clock_1_out_nativeaddress,
      master_read => nios2_clock_1_out_read,
      master_write => nios2_clock_1_out_write,
      master_writedata => nios2_clock_1_out_writedata,
      slave_endofpacket => nios2_clock_1_in_endofpacket,
      slave_readdata => nios2_clock_1_in_readdata,
      slave_waitrequest => nios2_clock_1_in_waitrequest,
      master_clk => internal_altpll_0_c0,
      master_endofpacket => nios2_clock_1_out_endofpacket,
      master_readdata => nios2_clock_1_out_readdata,
      master_reset_n => nios2_clock_1_out_reset_n,
      master_waitrequest => nios2_clock_1_out_waitrequest,
      slave_address => nios2_clock_1_in_address,
      slave_byteenable => nios2_clock_1_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_1_in_nativeaddress,
      slave_read => nios2_clock_1_in_read,
      slave_reset_n => nios2_clock_1_in_reset_n,
      slave_write => nios2_clock_1_in_write,
      slave_writedata => nios2_clock_1_in_writedata
    );


  --the_nios2_clock_10_in, which is an e_instance
  the_nios2_clock_10_in : nios2_clock_10_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_10_in => cpu_0_data_master_granted_nios2_clock_10_in,
      cpu_0_data_master_qualified_request_nios2_clock_10_in => cpu_0_data_master_qualified_request_nios2_clock_10_in,
      cpu_0_data_master_read_data_valid_nios2_clock_10_in => cpu_0_data_master_read_data_valid_nios2_clock_10_in,
      cpu_0_data_master_requests_nios2_clock_10_in => cpu_0_data_master_requests_nios2_clock_10_in,
      d1_nios2_clock_10_in_end_xfer => d1_nios2_clock_10_in_end_xfer,
      nios2_clock_10_in_address => nios2_clock_10_in_address,
      nios2_clock_10_in_endofpacket_from_sa => nios2_clock_10_in_endofpacket_from_sa,
      nios2_clock_10_in_nativeaddress => nios2_clock_10_in_nativeaddress,
      nios2_clock_10_in_read => nios2_clock_10_in_read,
      nios2_clock_10_in_readdata_from_sa => nios2_clock_10_in_readdata_from_sa,
      nios2_clock_10_in_reset_n => nios2_clock_10_in_reset_n,
      nios2_clock_10_in_waitrequest_from_sa => nios2_clock_10_in_waitrequest_from_sa,
      nios2_clock_10_in_write => nios2_clock_10_in_write,
      nios2_clock_10_in_writedata => nios2_clock_10_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_10_in_endofpacket => nios2_clock_10_in_endofpacket,
      nios2_clock_10_in_readdata => nios2_clock_10_in_readdata,
      nios2_clock_10_in_waitrequest => nios2_clock_10_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_10_out, which is an e_instance
  the_nios2_clock_10_out : nios2_clock_10_out_arbitrator
    port map(
      nios2_clock_10_out_address_to_slave => nios2_clock_10_out_address_to_slave,
      nios2_clock_10_out_readdata => nios2_clock_10_out_readdata,
      nios2_clock_10_out_reset_n => nios2_clock_10_out_reset_n,
      nios2_clock_10_out_waitrequest => nios2_clock_10_out_waitrequest,
      clk => internal_altpll_0_c0,
      d1_mode_select_s1_end_xfer => d1_mode_select_s1_end_xfer,
      mode_select_s1_readdata_from_sa => mode_select_s1_readdata_from_sa,
      nios2_clock_10_out_address => nios2_clock_10_out_address,
      nios2_clock_10_out_granted_mode_select_s1 => nios2_clock_10_out_granted_mode_select_s1,
      nios2_clock_10_out_qualified_request_mode_select_s1 => nios2_clock_10_out_qualified_request_mode_select_s1,
      nios2_clock_10_out_read => nios2_clock_10_out_read,
      nios2_clock_10_out_read_data_valid_mode_select_s1 => nios2_clock_10_out_read_data_valid_mode_select_s1,
      nios2_clock_10_out_requests_mode_select_s1 => nios2_clock_10_out_requests_mode_select_s1,
      nios2_clock_10_out_write => nios2_clock_10_out_write,
      nios2_clock_10_out_writedata => nios2_clock_10_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_nios2_clock_10, which is an e_ptf_instance
  the_nios2_clock_10 : nios2_clock_10
    port map(
      master_address => nios2_clock_10_out_address,
      master_nativeaddress => nios2_clock_10_out_nativeaddress,
      master_read => nios2_clock_10_out_read,
      master_write => nios2_clock_10_out_write,
      master_writedata => nios2_clock_10_out_writedata,
      slave_endofpacket => nios2_clock_10_in_endofpacket,
      slave_readdata => nios2_clock_10_in_readdata,
      slave_waitrequest => nios2_clock_10_in_waitrequest,
      master_clk => internal_altpll_0_c0,
      master_endofpacket => nios2_clock_10_out_endofpacket,
      master_readdata => nios2_clock_10_out_readdata,
      master_reset_n => nios2_clock_10_out_reset_n,
      master_waitrequest => nios2_clock_10_out_waitrequest,
      slave_address => nios2_clock_10_in_address,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_10_in_nativeaddress,
      slave_read => nios2_clock_10_in_read,
      slave_reset_n => nios2_clock_10_in_reset_n,
      slave_write => nios2_clock_10_in_write,
      slave_writedata => nios2_clock_10_in_writedata
    );


  --the_nios2_clock_11_in, which is an e_instance
  the_nios2_clock_11_in : nios2_clock_11_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_11_in => cpu_0_data_master_granted_nios2_clock_11_in,
      cpu_0_data_master_qualified_request_nios2_clock_11_in => cpu_0_data_master_qualified_request_nios2_clock_11_in,
      cpu_0_data_master_read_data_valid_nios2_clock_11_in => cpu_0_data_master_read_data_valid_nios2_clock_11_in,
      cpu_0_data_master_requests_nios2_clock_11_in => cpu_0_data_master_requests_nios2_clock_11_in,
      d1_nios2_clock_11_in_end_xfer => d1_nios2_clock_11_in_end_xfer,
      nios2_clock_11_in_address => nios2_clock_11_in_address,
      nios2_clock_11_in_endofpacket_from_sa => nios2_clock_11_in_endofpacket_from_sa,
      nios2_clock_11_in_nativeaddress => nios2_clock_11_in_nativeaddress,
      nios2_clock_11_in_read => nios2_clock_11_in_read,
      nios2_clock_11_in_readdata_from_sa => nios2_clock_11_in_readdata_from_sa,
      nios2_clock_11_in_reset_n => nios2_clock_11_in_reset_n,
      nios2_clock_11_in_waitrequest_from_sa => nios2_clock_11_in_waitrequest_from_sa,
      nios2_clock_11_in_write => nios2_clock_11_in_write,
      nios2_clock_11_in_writedata => nios2_clock_11_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_11_in_endofpacket => nios2_clock_11_in_endofpacket,
      nios2_clock_11_in_readdata => nios2_clock_11_in_readdata,
      nios2_clock_11_in_waitrequest => nios2_clock_11_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_11_out, which is an e_instance
  the_nios2_clock_11_out : nios2_clock_11_out_arbitrator
    port map(
      nios2_clock_11_out_address_to_slave => nios2_clock_11_out_address_to_slave,
      nios2_clock_11_out_readdata => nios2_clock_11_out_readdata,
      nios2_clock_11_out_reset_n => nios2_clock_11_out_reset_n,
      nios2_clock_11_out_waitrequest => nios2_clock_11_out_waitrequest,
      clk => internal_altpll_0_c0,
      comparator_pio_s1_readdata_from_sa => comparator_pio_s1_readdata_from_sa,
      d1_comparator_pio_s1_end_xfer => d1_comparator_pio_s1_end_xfer,
      nios2_clock_11_out_address => nios2_clock_11_out_address,
      nios2_clock_11_out_granted_comparator_pio_s1 => nios2_clock_11_out_granted_comparator_pio_s1,
      nios2_clock_11_out_qualified_request_comparator_pio_s1 => nios2_clock_11_out_qualified_request_comparator_pio_s1,
      nios2_clock_11_out_read => nios2_clock_11_out_read,
      nios2_clock_11_out_read_data_valid_comparator_pio_s1 => nios2_clock_11_out_read_data_valid_comparator_pio_s1,
      nios2_clock_11_out_requests_comparator_pio_s1 => nios2_clock_11_out_requests_comparator_pio_s1,
      nios2_clock_11_out_write => nios2_clock_11_out_write,
      nios2_clock_11_out_writedata => nios2_clock_11_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_nios2_clock_11, which is an e_ptf_instance
  the_nios2_clock_11 : nios2_clock_11
    port map(
      master_address => nios2_clock_11_out_address,
      master_nativeaddress => nios2_clock_11_out_nativeaddress,
      master_read => nios2_clock_11_out_read,
      master_write => nios2_clock_11_out_write,
      master_writedata => nios2_clock_11_out_writedata,
      slave_endofpacket => nios2_clock_11_in_endofpacket,
      slave_readdata => nios2_clock_11_in_readdata,
      slave_waitrequest => nios2_clock_11_in_waitrequest,
      master_clk => internal_altpll_0_c0,
      master_endofpacket => nios2_clock_11_out_endofpacket,
      master_readdata => nios2_clock_11_out_readdata,
      master_reset_n => nios2_clock_11_out_reset_n,
      master_waitrequest => nios2_clock_11_out_waitrequest,
      slave_address => nios2_clock_11_in_address,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_11_in_nativeaddress,
      slave_read => nios2_clock_11_in_read,
      slave_reset_n => nios2_clock_11_in_reset_n,
      slave_write => nios2_clock_11_in_write,
      slave_writedata => nios2_clock_11_in_writedata
    );


  --the_nios2_clock_12_in, which is an e_instance
  the_nios2_clock_12_in : nios2_clock_12_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_12_in => cpu_0_data_master_granted_nios2_clock_12_in,
      cpu_0_data_master_qualified_request_nios2_clock_12_in => cpu_0_data_master_qualified_request_nios2_clock_12_in,
      cpu_0_data_master_read_data_valid_nios2_clock_12_in => cpu_0_data_master_read_data_valid_nios2_clock_12_in,
      cpu_0_data_master_requests_nios2_clock_12_in => cpu_0_data_master_requests_nios2_clock_12_in,
      d1_nios2_clock_12_in_end_xfer => d1_nios2_clock_12_in_end_xfer,
      nios2_clock_12_in_address => nios2_clock_12_in_address,
      nios2_clock_12_in_endofpacket_from_sa => nios2_clock_12_in_endofpacket_from_sa,
      nios2_clock_12_in_nativeaddress => nios2_clock_12_in_nativeaddress,
      nios2_clock_12_in_read => nios2_clock_12_in_read,
      nios2_clock_12_in_readdata_from_sa => nios2_clock_12_in_readdata_from_sa,
      nios2_clock_12_in_reset_n => nios2_clock_12_in_reset_n,
      nios2_clock_12_in_waitrequest_from_sa => nios2_clock_12_in_waitrequest_from_sa,
      nios2_clock_12_in_write => nios2_clock_12_in_write,
      nios2_clock_12_in_writedata => nios2_clock_12_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_12_in_endofpacket => nios2_clock_12_in_endofpacket,
      nios2_clock_12_in_readdata => nios2_clock_12_in_readdata,
      nios2_clock_12_in_waitrequest => nios2_clock_12_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_12_out, which is an e_instance
  the_nios2_clock_12_out : nios2_clock_12_out_arbitrator
    port map(
      nios2_clock_12_out_address_to_slave => nios2_clock_12_out_address_to_slave,
      nios2_clock_12_out_readdata => nios2_clock_12_out_readdata,
      nios2_clock_12_out_reset_n => nios2_clock_12_out_reset_n,
      nios2_clock_12_out_waitrequest => nios2_clock_12_out_waitrequest,
      clk => clk_0,
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      nios2_clock_12_out_address => nios2_clock_12_out_address,
      nios2_clock_12_out_granted_led_pio_s1 => nios2_clock_12_out_granted_led_pio_s1,
      nios2_clock_12_out_qualified_request_led_pio_s1 => nios2_clock_12_out_qualified_request_led_pio_s1,
      nios2_clock_12_out_read => nios2_clock_12_out_read,
      nios2_clock_12_out_read_data_valid_led_pio_s1 => nios2_clock_12_out_read_data_valid_led_pio_s1,
      nios2_clock_12_out_requests_led_pio_s1 => nios2_clock_12_out_requests_led_pio_s1,
      nios2_clock_12_out_write => nios2_clock_12_out_write,
      nios2_clock_12_out_writedata => nios2_clock_12_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_nios2_clock_12, which is an e_ptf_instance
  the_nios2_clock_12 : nios2_clock_12
    port map(
      master_address => nios2_clock_12_out_address,
      master_nativeaddress => nios2_clock_12_out_nativeaddress,
      master_read => nios2_clock_12_out_read,
      master_write => nios2_clock_12_out_write,
      master_writedata => nios2_clock_12_out_writedata,
      slave_endofpacket => nios2_clock_12_in_endofpacket,
      slave_readdata => nios2_clock_12_in_readdata,
      slave_waitrequest => nios2_clock_12_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_12_out_endofpacket,
      master_readdata => nios2_clock_12_out_readdata,
      master_reset_n => nios2_clock_12_out_reset_n,
      master_waitrequest => nios2_clock_12_out_waitrequest,
      slave_address => nios2_clock_12_in_address,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_12_in_nativeaddress,
      slave_read => nios2_clock_12_in_read,
      slave_reset_n => nios2_clock_12_in_reset_n,
      slave_write => nios2_clock_12_in_write,
      slave_writedata => nios2_clock_12_in_writedata
    );


  --the_nios2_clock_13_in, which is an e_instance
  the_nios2_clock_13_in : nios2_clock_13_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_13_in => cpu_0_data_master_granted_nios2_clock_13_in,
      cpu_0_data_master_qualified_request_nios2_clock_13_in => cpu_0_data_master_qualified_request_nios2_clock_13_in,
      cpu_0_data_master_read_data_valid_nios2_clock_13_in => cpu_0_data_master_read_data_valid_nios2_clock_13_in,
      cpu_0_data_master_requests_nios2_clock_13_in => cpu_0_data_master_requests_nios2_clock_13_in,
      d1_nios2_clock_13_in_end_xfer => d1_nios2_clock_13_in_end_xfer,
      nios2_clock_13_in_address => nios2_clock_13_in_address,
      nios2_clock_13_in_endofpacket_from_sa => nios2_clock_13_in_endofpacket_from_sa,
      nios2_clock_13_in_nativeaddress => nios2_clock_13_in_nativeaddress,
      nios2_clock_13_in_read => nios2_clock_13_in_read,
      nios2_clock_13_in_readdata_from_sa => nios2_clock_13_in_readdata_from_sa,
      nios2_clock_13_in_reset_n => nios2_clock_13_in_reset_n,
      nios2_clock_13_in_waitrequest_from_sa => nios2_clock_13_in_waitrequest_from_sa,
      nios2_clock_13_in_write => nios2_clock_13_in_write,
      nios2_clock_13_in_writedata => nios2_clock_13_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_13_in_endofpacket => nios2_clock_13_in_endofpacket,
      nios2_clock_13_in_readdata => nios2_clock_13_in_readdata,
      nios2_clock_13_in_waitrequest => nios2_clock_13_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_13_out, which is an e_instance
  the_nios2_clock_13_out : nios2_clock_13_out_arbitrator
    port map(
      nios2_clock_13_out_address_to_slave => nios2_clock_13_out_address_to_slave,
      nios2_clock_13_out_readdata => nios2_clock_13_out_readdata,
      nios2_clock_13_out_reset_n => nios2_clock_13_out_reset_n,
      nios2_clock_13_out_waitrequest => nios2_clock_13_out_waitrequest,
      clk => clk_0,
      d1_gen_code_strobe_s1_end_xfer => d1_gen_code_strobe_s1_end_xfer,
      gen_code_strobe_s1_readdata_from_sa => gen_code_strobe_s1_readdata_from_sa,
      nios2_clock_13_out_address => nios2_clock_13_out_address,
      nios2_clock_13_out_granted_gen_code_strobe_s1 => nios2_clock_13_out_granted_gen_code_strobe_s1,
      nios2_clock_13_out_qualified_request_gen_code_strobe_s1 => nios2_clock_13_out_qualified_request_gen_code_strobe_s1,
      nios2_clock_13_out_read => nios2_clock_13_out_read,
      nios2_clock_13_out_read_data_valid_gen_code_strobe_s1 => nios2_clock_13_out_read_data_valid_gen_code_strobe_s1,
      nios2_clock_13_out_requests_gen_code_strobe_s1 => nios2_clock_13_out_requests_gen_code_strobe_s1,
      nios2_clock_13_out_write => nios2_clock_13_out_write,
      nios2_clock_13_out_writedata => nios2_clock_13_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_nios2_clock_13, which is an e_ptf_instance
  the_nios2_clock_13 : nios2_clock_13
    port map(
      master_address => nios2_clock_13_out_address,
      master_nativeaddress => nios2_clock_13_out_nativeaddress,
      master_read => nios2_clock_13_out_read,
      master_write => nios2_clock_13_out_write,
      master_writedata => nios2_clock_13_out_writedata,
      slave_endofpacket => nios2_clock_13_in_endofpacket,
      slave_readdata => nios2_clock_13_in_readdata,
      slave_waitrequest => nios2_clock_13_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_13_out_endofpacket,
      master_readdata => nios2_clock_13_out_readdata,
      master_reset_n => nios2_clock_13_out_reset_n,
      master_waitrequest => nios2_clock_13_out_waitrequest,
      slave_address => nios2_clock_13_in_address,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_13_in_nativeaddress,
      slave_read => nios2_clock_13_in_read,
      slave_reset_n => nios2_clock_13_in_reset_n,
      slave_write => nios2_clock_13_in_write,
      slave_writedata => nios2_clock_13_in_writedata
    );


  --the_nios2_clock_14_in, which is an e_instance
  the_nios2_clock_14_in : nios2_clock_14_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_14_in => cpu_0_data_master_granted_nios2_clock_14_in,
      cpu_0_data_master_qualified_request_nios2_clock_14_in => cpu_0_data_master_qualified_request_nios2_clock_14_in,
      cpu_0_data_master_read_data_valid_nios2_clock_14_in => cpu_0_data_master_read_data_valid_nios2_clock_14_in,
      cpu_0_data_master_requests_nios2_clock_14_in => cpu_0_data_master_requests_nios2_clock_14_in,
      d1_nios2_clock_14_in_end_xfer => d1_nios2_clock_14_in_end_xfer,
      nios2_clock_14_in_address => nios2_clock_14_in_address,
      nios2_clock_14_in_endofpacket_from_sa => nios2_clock_14_in_endofpacket_from_sa,
      nios2_clock_14_in_nativeaddress => nios2_clock_14_in_nativeaddress,
      nios2_clock_14_in_read => nios2_clock_14_in_read,
      nios2_clock_14_in_readdata_from_sa => nios2_clock_14_in_readdata_from_sa,
      nios2_clock_14_in_reset_n => nios2_clock_14_in_reset_n,
      nios2_clock_14_in_waitrequest_from_sa => nios2_clock_14_in_waitrequest_from_sa,
      nios2_clock_14_in_write => nios2_clock_14_in_write,
      nios2_clock_14_in_writedata => nios2_clock_14_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_14_in_endofpacket => nios2_clock_14_in_endofpacket,
      nios2_clock_14_in_readdata => nios2_clock_14_in_readdata,
      nios2_clock_14_in_waitrequest => nios2_clock_14_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_14_out, which is an e_instance
  the_nios2_clock_14_out : nios2_clock_14_out_arbitrator
    port map(
      nios2_clock_14_out_address_to_slave => nios2_clock_14_out_address_to_slave,
      nios2_clock_14_out_readdata => nios2_clock_14_out_readdata,
      nios2_clock_14_out_reset_n => nios2_clock_14_out_reset_n,
      nios2_clock_14_out_waitrequest => nios2_clock_14_out_waitrequest,
      clk => clk_0,
      d1_switch_pio_s1_end_xfer => d1_switch_pio_s1_end_xfer,
      nios2_clock_14_out_address => nios2_clock_14_out_address,
      nios2_clock_14_out_granted_switch_pio_s1 => nios2_clock_14_out_granted_switch_pio_s1,
      nios2_clock_14_out_qualified_request_switch_pio_s1 => nios2_clock_14_out_qualified_request_switch_pio_s1,
      nios2_clock_14_out_read => nios2_clock_14_out_read,
      nios2_clock_14_out_read_data_valid_switch_pio_s1 => nios2_clock_14_out_read_data_valid_switch_pio_s1,
      nios2_clock_14_out_requests_switch_pio_s1 => nios2_clock_14_out_requests_switch_pio_s1,
      nios2_clock_14_out_write => nios2_clock_14_out_write,
      nios2_clock_14_out_writedata => nios2_clock_14_out_writedata,
      reset_n => clk_0_reset_n,
      switch_pio_s1_readdata_from_sa => switch_pio_s1_readdata_from_sa
    );


  --the_nios2_clock_14, which is an e_ptf_instance
  the_nios2_clock_14 : nios2_clock_14
    port map(
      master_address => nios2_clock_14_out_address,
      master_nativeaddress => nios2_clock_14_out_nativeaddress,
      master_read => nios2_clock_14_out_read,
      master_write => nios2_clock_14_out_write,
      master_writedata => nios2_clock_14_out_writedata,
      slave_endofpacket => nios2_clock_14_in_endofpacket,
      slave_readdata => nios2_clock_14_in_readdata,
      slave_waitrequest => nios2_clock_14_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_14_out_endofpacket,
      master_readdata => nios2_clock_14_out_readdata,
      master_reset_n => nios2_clock_14_out_reset_n,
      master_waitrequest => nios2_clock_14_out_waitrequest,
      slave_address => nios2_clock_14_in_address,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_14_in_nativeaddress,
      slave_read => nios2_clock_14_in_read,
      slave_reset_n => nios2_clock_14_in_reset_n,
      slave_write => nios2_clock_14_in_write,
      slave_writedata => nios2_clock_14_in_writedata
    );


  --the_nios2_clock_15_in, which is an e_instance
  the_nios2_clock_15_in : nios2_clock_15_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_15_in => cpu_0_data_master_granted_nios2_clock_15_in,
      cpu_0_data_master_qualified_request_nios2_clock_15_in => cpu_0_data_master_qualified_request_nios2_clock_15_in,
      cpu_0_data_master_read_data_valid_nios2_clock_15_in => cpu_0_data_master_read_data_valid_nios2_clock_15_in,
      cpu_0_data_master_requests_nios2_clock_15_in => cpu_0_data_master_requests_nios2_clock_15_in,
      d1_nios2_clock_15_in_end_xfer => d1_nios2_clock_15_in_end_xfer,
      nios2_clock_15_in_address => nios2_clock_15_in_address,
      nios2_clock_15_in_byteenable => nios2_clock_15_in_byteenable,
      nios2_clock_15_in_endofpacket_from_sa => nios2_clock_15_in_endofpacket_from_sa,
      nios2_clock_15_in_nativeaddress => nios2_clock_15_in_nativeaddress,
      nios2_clock_15_in_read => nios2_clock_15_in_read,
      nios2_clock_15_in_readdata_from_sa => nios2_clock_15_in_readdata_from_sa,
      nios2_clock_15_in_reset_n => nios2_clock_15_in_reset_n,
      nios2_clock_15_in_waitrequest_from_sa => nios2_clock_15_in_waitrequest_from_sa,
      nios2_clock_15_in_write => nios2_clock_15_in_write,
      nios2_clock_15_in_writedata => nios2_clock_15_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_15_in_endofpacket => nios2_clock_15_in_endofpacket,
      nios2_clock_15_in_readdata => nios2_clock_15_in_readdata,
      nios2_clock_15_in_waitrequest => nios2_clock_15_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_15_out, which is an e_instance
  the_nios2_clock_15_out : nios2_clock_15_out_arbitrator
    port map(
      nios2_clock_15_out_address_to_slave => nios2_clock_15_out_address_to_slave,
      nios2_clock_15_out_readdata => nios2_clock_15_out_readdata,
      nios2_clock_15_out_reset_n => nios2_clock_15_out_reset_n,
      nios2_clock_15_out_waitrequest => nios2_clock_15_out_waitrequest,
      cal_dac_code_pio_s1_readdata_from_sa => cal_dac_code_pio_s1_readdata_from_sa,
      clk => clk_0,
      d1_cal_dac_code_pio_s1_end_xfer => d1_cal_dac_code_pio_s1_end_xfer,
      nios2_clock_15_out_address => nios2_clock_15_out_address,
      nios2_clock_15_out_byteenable => nios2_clock_15_out_byteenable,
      nios2_clock_15_out_granted_cal_dac_code_pio_s1 => nios2_clock_15_out_granted_cal_dac_code_pio_s1,
      nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1 => nios2_clock_15_out_qualified_request_cal_dac_code_pio_s1,
      nios2_clock_15_out_read => nios2_clock_15_out_read,
      nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1 => nios2_clock_15_out_read_data_valid_cal_dac_code_pio_s1,
      nios2_clock_15_out_requests_cal_dac_code_pio_s1 => nios2_clock_15_out_requests_cal_dac_code_pio_s1,
      nios2_clock_15_out_write => nios2_clock_15_out_write,
      nios2_clock_15_out_writedata => nios2_clock_15_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_nios2_clock_15, which is an e_ptf_instance
  the_nios2_clock_15 : nios2_clock_15
    port map(
      master_address => nios2_clock_15_out_address,
      master_byteenable => nios2_clock_15_out_byteenable,
      master_nativeaddress => nios2_clock_15_out_nativeaddress,
      master_read => nios2_clock_15_out_read,
      master_write => nios2_clock_15_out_write,
      master_writedata => nios2_clock_15_out_writedata,
      slave_endofpacket => nios2_clock_15_in_endofpacket,
      slave_readdata => nios2_clock_15_in_readdata,
      slave_waitrequest => nios2_clock_15_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_15_out_endofpacket,
      master_readdata => nios2_clock_15_out_readdata,
      master_reset_n => nios2_clock_15_out_reset_n,
      master_waitrequest => nios2_clock_15_out_waitrequest,
      slave_address => nios2_clock_15_in_address,
      slave_byteenable => nios2_clock_15_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_15_in_nativeaddress,
      slave_read => nios2_clock_15_in_read,
      slave_reset_n => nios2_clock_15_in_reset_n,
      slave_write => nios2_clock_15_in_write,
      slave_writedata => nios2_clock_15_in_writedata
    );


  --the_nios2_clock_16_in, which is an e_instance
  the_nios2_clock_16_in : nios2_clock_16_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_16_in => cpu_0_data_master_granted_nios2_clock_16_in,
      cpu_0_data_master_qualified_request_nios2_clock_16_in => cpu_0_data_master_qualified_request_nios2_clock_16_in,
      cpu_0_data_master_read_data_valid_nios2_clock_16_in => cpu_0_data_master_read_data_valid_nios2_clock_16_in,
      cpu_0_data_master_requests_nios2_clock_16_in => cpu_0_data_master_requests_nios2_clock_16_in,
      d1_nios2_clock_16_in_end_xfer => d1_nios2_clock_16_in_end_xfer,
      nios2_clock_16_in_address => nios2_clock_16_in_address,
      nios2_clock_16_in_byteenable => nios2_clock_16_in_byteenable,
      nios2_clock_16_in_endofpacket_from_sa => nios2_clock_16_in_endofpacket_from_sa,
      nios2_clock_16_in_nativeaddress => nios2_clock_16_in_nativeaddress,
      nios2_clock_16_in_read => nios2_clock_16_in_read,
      nios2_clock_16_in_readdata_from_sa => nios2_clock_16_in_readdata_from_sa,
      nios2_clock_16_in_reset_n => nios2_clock_16_in_reset_n,
      nios2_clock_16_in_waitrequest_from_sa => nios2_clock_16_in_waitrequest_from_sa,
      nios2_clock_16_in_write => nios2_clock_16_in_write,
      nios2_clock_16_in_writedata => nios2_clock_16_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_16_in_endofpacket => nios2_clock_16_in_endofpacket,
      nios2_clock_16_in_readdata => nios2_clock_16_in_readdata,
      nios2_clock_16_in_waitrequest => nios2_clock_16_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_16_out, which is an e_instance
  the_nios2_clock_16_out : nios2_clock_16_out_arbitrator
    port map(
      nios2_clock_16_out_address_to_slave => nios2_clock_16_out_address_to_slave,
      nios2_clock_16_out_readdata => nios2_clock_16_out_readdata,
      nios2_clock_16_out_reset_n => nios2_clock_16_out_reset_n,
      nios2_clock_16_out_waitrequest => nios2_clock_16_out_waitrequest,
      clk => clk_0,
      d1_usb_code_pio_s1_end_xfer => d1_usb_code_pio_s1_end_xfer,
      nios2_clock_16_out_address => nios2_clock_16_out_address,
      nios2_clock_16_out_byteenable => nios2_clock_16_out_byteenable,
      nios2_clock_16_out_granted_usb_code_pio_s1 => nios2_clock_16_out_granted_usb_code_pio_s1,
      nios2_clock_16_out_qualified_request_usb_code_pio_s1 => nios2_clock_16_out_qualified_request_usb_code_pio_s1,
      nios2_clock_16_out_read => nios2_clock_16_out_read,
      nios2_clock_16_out_read_data_valid_usb_code_pio_s1 => nios2_clock_16_out_read_data_valid_usb_code_pio_s1,
      nios2_clock_16_out_requests_usb_code_pio_s1 => nios2_clock_16_out_requests_usb_code_pio_s1,
      nios2_clock_16_out_write => nios2_clock_16_out_write,
      nios2_clock_16_out_writedata => nios2_clock_16_out_writedata,
      reset_n => clk_0_reset_n,
      usb_code_pio_s1_readdata_from_sa => usb_code_pio_s1_readdata_from_sa
    );


  --the_nios2_clock_16, which is an e_ptf_instance
  the_nios2_clock_16 : nios2_clock_16
    port map(
      master_address => nios2_clock_16_out_address,
      master_byteenable => nios2_clock_16_out_byteenable,
      master_nativeaddress => nios2_clock_16_out_nativeaddress,
      master_read => nios2_clock_16_out_read,
      master_write => nios2_clock_16_out_write,
      master_writedata => nios2_clock_16_out_writedata,
      slave_endofpacket => nios2_clock_16_in_endofpacket,
      slave_readdata => nios2_clock_16_in_readdata,
      slave_waitrequest => nios2_clock_16_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_16_out_endofpacket,
      master_readdata => nios2_clock_16_out_readdata,
      master_reset_n => nios2_clock_16_out_reset_n,
      master_waitrequest => nios2_clock_16_out_waitrequest,
      slave_address => nios2_clock_16_in_address,
      slave_byteenable => nios2_clock_16_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_16_in_nativeaddress,
      slave_read => nios2_clock_16_in_read,
      slave_reset_n => nios2_clock_16_in_reset_n,
      slave_write => nios2_clock_16_in_write,
      slave_writedata => nios2_clock_16_in_writedata
    );


  --the_nios2_clock_17_in, which is an e_instance
  the_nios2_clock_17_in : nios2_clock_17_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_17_in => cpu_0_data_master_granted_nios2_clock_17_in,
      cpu_0_data_master_qualified_request_nios2_clock_17_in => cpu_0_data_master_qualified_request_nios2_clock_17_in,
      cpu_0_data_master_read_data_valid_nios2_clock_17_in => cpu_0_data_master_read_data_valid_nios2_clock_17_in,
      cpu_0_data_master_requests_nios2_clock_17_in => cpu_0_data_master_requests_nios2_clock_17_in,
      d1_nios2_clock_17_in_end_xfer => d1_nios2_clock_17_in_end_xfer,
      nios2_clock_17_in_address => nios2_clock_17_in_address,
      nios2_clock_17_in_endofpacket_from_sa => nios2_clock_17_in_endofpacket_from_sa,
      nios2_clock_17_in_nativeaddress => nios2_clock_17_in_nativeaddress,
      nios2_clock_17_in_read => nios2_clock_17_in_read,
      nios2_clock_17_in_readdata_from_sa => nios2_clock_17_in_readdata_from_sa,
      nios2_clock_17_in_reset_n => nios2_clock_17_in_reset_n,
      nios2_clock_17_in_waitrequest_from_sa => nios2_clock_17_in_waitrequest_from_sa,
      nios2_clock_17_in_write => nios2_clock_17_in_write,
      nios2_clock_17_in_writedata => nios2_clock_17_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_17_in_endofpacket => nios2_clock_17_in_endofpacket,
      nios2_clock_17_in_readdata => nios2_clock_17_in_readdata,
      nios2_clock_17_in_waitrequest => nios2_clock_17_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_17_out, which is an e_instance
  the_nios2_clock_17_out : nios2_clock_17_out_arbitrator
    port map(
      nios2_clock_17_out_address_to_slave => nios2_clock_17_out_address_to_slave,
      nios2_clock_17_out_readdata => nios2_clock_17_out_readdata,
      nios2_clock_17_out_reset_n => nios2_clock_17_out_reset_n,
      nios2_clock_17_out_waitrequest => nios2_clock_17_out_waitrequest,
      clk => clk_0,
      d1_sample_and_hold_pio_s1_end_xfer => d1_sample_and_hold_pio_s1_end_xfer,
      nios2_clock_17_out_address => nios2_clock_17_out_address,
      nios2_clock_17_out_granted_sample_and_hold_pio_s1 => nios2_clock_17_out_granted_sample_and_hold_pio_s1,
      nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 => nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1,
      nios2_clock_17_out_read => nios2_clock_17_out_read,
      nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1 => nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1,
      nios2_clock_17_out_requests_sample_and_hold_pio_s1 => nios2_clock_17_out_requests_sample_and_hold_pio_s1,
      nios2_clock_17_out_write => nios2_clock_17_out_write,
      nios2_clock_17_out_writedata => nios2_clock_17_out_writedata,
      reset_n => clk_0_reset_n,
      sample_and_hold_pio_s1_readdata_from_sa => sample_and_hold_pio_s1_readdata_from_sa
    );


  --the_nios2_clock_17, which is an e_ptf_instance
  the_nios2_clock_17 : nios2_clock_17
    port map(
      master_address => nios2_clock_17_out_address,
      master_nativeaddress => nios2_clock_17_out_nativeaddress,
      master_read => nios2_clock_17_out_read,
      master_write => nios2_clock_17_out_write,
      master_writedata => nios2_clock_17_out_writedata,
      slave_endofpacket => nios2_clock_17_in_endofpacket,
      slave_readdata => nios2_clock_17_in_readdata,
      slave_waitrequest => nios2_clock_17_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_17_out_endofpacket,
      master_readdata => nios2_clock_17_out_readdata,
      master_reset_n => nios2_clock_17_out_reset_n,
      master_waitrequest => nios2_clock_17_out_waitrequest,
      slave_address => nios2_clock_17_in_address,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_17_in_nativeaddress,
      slave_read => nios2_clock_17_in_read,
      slave_reset_n => nios2_clock_17_in_reset_n,
      slave_write => nios2_clock_17_in_write,
      slave_writedata => nios2_clock_17_in_writedata
    );


  --the_nios2_clock_18_in, which is an e_instance
  the_nios2_clock_18_in : nios2_clock_18_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_18_in => cpu_0_data_master_granted_nios2_clock_18_in,
      cpu_0_data_master_qualified_request_nios2_clock_18_in => cpu_0_data_master_qualified_request_nios2_clock_18_in,
      cpu_0_data_master_read_data_valid_nios2_clock_18_in => cpu_0_data_master_read_data_valid_nios2_clock_18_in,
      cpu_0_data_master_requests_nios2_clock_18_in => cpu_0_data_master_requests_nios2_clock_18_in,
      d1_nios2_clock_18_in_end_xfer => d1_nios2_clock_18_in_end_xfer,
      nios2_clock_18_in_address => nios2_clock_18_in_address,
      nios2_clock_18_in_endofpacket_from_sa => nios2_clock_18_in_endofpacket_from_sa,
      nios2_clock_18_in_nativeaddress => nios2_clock_18_in_nativeaddress,
      nios2_clock_18_in_read => nios2_clock_18_in_read,
      nios2_clock_18_in_readdata_from_sa => nios2_clock_18_in_readdata_from_sa,
      nios2_clock_18_in_reset_n => nios2_clock_18_in_reset_n,
      nios2_clock_18_in_waitrequest_from_sa => nios2_clock_18_in_waitrequest_from_sa,
      nios2_clock_18_in_write => nios2_clock_18_in_write,
      nios2_clock_18_in_writedata => nios2_clock_18_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_18_in_endofpacket => nios2_clock_18_in_endofpacket,
      nios2_clock_18_in_readdata => nios2_clock_18_in_readdata,
      nios2_clock_18_in_waitrequest => nios2_clock_18_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_18_out, which is an e_instance
  the_nios2_clock_18_out : nios2_clock_18_out_arbitrator
    port map(
      nios2_clock_18_out_address_to_slave => nios2_clock_18_out_address_to_slave,
      nios2_clock_18_out_readdata => nios2_clock_18_out_readdata,
      nios2_clock_18_out_reset_n => nios2_clock_18_out_reset_n,
      nios2_clock_18_out_waitrequest => nios2_clock_18_out_waitrequest,
      clk => clk_0,
      d1_latch_pio_s1_end_xfer => d1_latch_pio_s1_end_xfer,
      latch_pio_s1_readdata_from_sa => latch_pio_s1_readdata_from_sa,
      nios2_clock_18_out_address => nios2_clock_18_out_address,
      nios2_clock_18_out_granted_latch_pio_s1 => nios2_clock_18_out_granted_latch_pio_s1,
      nios2_clock_18_out_qualified_request_latch_pio_s1 => nios2_clock_18_out_qualified_request_latch_pio_s1,
      nios2_clock_18_out_read => nios2_clock_18_out_read,
      nios2_clock_18_out_read_data_valid_latch_pio_s1 => nios2_clock_18_out_read_data_valid_latch_pio_s1,
      nios2_clock_18_out_requests_latch_pio_s1 => nios2_clock_18_out_requests_latch_pio_s1,
      nios2_clock_18_out_write => nios2_clock_18_out_write,
      nios2_clock_18_out_writedata => nios2_clock_18_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_nios2_clock_18, which is an e_ptf_instance
  the_nios2_clock_18 : nios2_clock_18
    port map(
      master_address => nios2_clock_18_out_address,
      master_nativeaddress => nios2_clock_18_out_nativeaddress,
      master_read => nios2_clock_18_out_read,
      master_write => nios2_clock_18_out_write,
      master_writedata => nios2_clock_18_out_writedata,
      slave_endofpacket => nios2_clock_18_in_endofpacket,
      slave_readdata => nios2_clock_18_in_readdata,
      slave_waitrequest => nios2_clock_18_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_18_out_endofpacket,
      master_readdata => nios2_clock_18_out_readdata,
      master_reset_n => nios2_clock_18_out_reset_n,
      master_waitrequest => nios2_clock_18_out_waitrequest,
      slave_address => nios2_clock_18_in_address,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_18_in_nativeaddress,
      slave_read => nios2_clock_18_in_read,
      slave_reset_n => nios2_clock_18_in_reset_n,
      slave_write => nios2_clock_18_in_write,
      slave_writedata => nios2_clock_18_in_writedata
    );


  --the_nios2_clock_2_in, which is an e_instance
  the_nios2_clock_2_in : nios2_clock_2_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_2_in => cpu_0_data_master_granted_nios2_clock_2_in,
      cpu_0_data_master_qualified_request_nios2_clock_2_in => cpu_0_data_master_qualified_request_nios2_clock_2_in,
      cpu_0_data_master_read_data_valid_nios2_clock_2_in => cpu_0_data_master_read_data_valid_nios2_clock_2_in,
      cpu_0_data_master_requests_nios2_clock_2_in => cpu_0_data_master_requests_nios2_clock_2_in,
      d1_nios2_clock_2_in_end_xfer => d1_nios2_clock_2_in_end_xfer,
      nios2_clock_2_in_address => nios2_clock_2_in_address,
      nios2_clock_2_in_byteenable => nios2_clock_2_in_byteenable,
      nios2_clock_2_in_endofpacket_from_sa => nios2_clock_2_in_endofpacket_from_sa,
      nios2_clock_2_in_nativeaddress => nios2_clock_2_in_nativeaddress,
      nios2_clock_2_in_read => nios2_clock_2_in_read,
      nios2_clock_2_in_readdata_from_sa => nios2_clock_2_in_readdata_from_sa,
      nios2_clock_2_in_reset_n => nios2_clock_2_in_reset_n,
      nios2_clock_2_in_waitrequest_from_sa => nios2_clock_2_in_waitrequest_from_sa,
      nios2_clock_2_in_write => nios2_clock_2_in_write,
      nios2_clock_2_in_writedata => nios2_clock_2_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_2_in_endofpacket => nios2_clock_2_in_endofpacket,
      nios2_clock_2_in_readdata => nios2_clock_2_in_readdata,
      nios2_clock_2_in_waitrequest => nios2_clock_2_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_2_out, which is an e_instance
  the_nios2_clock_2_out : nios2_clock_2_out_arbitrator
    port map(
      nios2_clock_2_out_address_to_slave => nios2_clock_2_out_address_to_slave,
      nios2_clock_2_out_readdata => nios2_clock_2_out_readdata,
      nios2_clock_2_out_reset_n => nios2_clock_2_out_reset_n,
      nios2_clock_2_out_waitrequest => nios2_clock_2_out_waitrequest,
      clk => internal_altpll_0_c0,
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer => d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
      jtag_uart_0_avalon_jtag_slave_readdata_from_sa => jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
      nios2_clock_2_out_address => nios2_clock_2_out_address,
      nios2_clock_2_out_byteenable => nios2_clock_2_out_byteenable,
      nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_granted_jtag_uart_0_avalon_jtag_slave,
      nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_qualified_request_jtag_uart_0_avalon_jtag_slave,
      nios2_clock_2_out_read => nios2_clock_2_out_read,
      nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_read_data_valid_jtag_uart_0_avalon_jtag_slave,
      nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave => nios2_clock_2_out_requests_jtag_uart_0_avalon_jtag_slave,
      nios2_clock_2_out_write => nios2_clock_2_out_write,
      nios2_clock_2_out_writedata => nios2_clock_2_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_nios2_clock_2, which is an e_ptf_instance
  the_nios2_clock_2 : nios2_clock_2
    port map(
      master_address => nios2_clock_2_out_address,
      master_byteenable => nios2_clock_2_out_byteenable,
      master_nativeaddress => nios2_clock_2_out_nativeaddress,
      master_read => nios2_clock_2_out_read,
      master_write => nios2_clock_2_out_write,
      master_writedata => nios2_clock_2_out_writedata,
      slave_endofpacket => nios2_clock_2_in_endofpacket,
      slave_readdata => nios2_clock_2_in_readdata,
      slave_waitrequest => nios2_clock_2_in_waitrequest,
      master_clk => internal_altpll_0_c0,
      master_endofpacket => nios2_clock_2_out_endofpacket,
      master_readdata => nios2_clock_2_out_readdata,
      master_reset_n => nios2_clock_2_out_reset_n,
      master_waitrequest => nios2_clock_2_out_waitrequest,
      slave_address => nios2_clock_2_in_address,
      slave_byteenable => nios2_clock_2_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_2_in_nativeaddress,
      slave_read => nios2_clock_2_in_read,
      slave_reset_n => nios2_clock_2_in_reset_n,
      slave_write => nios2_clock_2_in_write,
      slave_writedata => nios2_clock_2_in_writedata
    );


  --the_nios2_clock_3_in, which is an e_instance
  the_nios2_clock_3_in : nios2_clock_3_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_3_in => cpu_0_data_master_granted_nios2_clock_3_in,
      cpu_0_data_master_qualified_request_nios2_clock_3_in => cpu_0_data_master_qualified_request_nios2_clock_3_in,
      cpu_0_data_master_read_data_valid_nios2_clock_3_in => cpu_0_data_master_read_data_valid_nios2_clock_3_in,
      cpu_0_data_master_requests_nios2_clock_3_in => cpu_0_data_master_requests_nios2_clock_3_in,
      d1_nios2_clock_3_in_end_xfer => d1_nios2_clock_3_in_end_xfer,
      nios2_clock_3_in_address => nios2_clock_3_in_address,
      nios2_clock_3_in_byteenable => nios2_clock_3_in_byteenable,
      nios2_clock_3_in_endofpacket_from_sa => nios2_clock_3_in_endofpacket_from_sa,
      nios2_clock_3_in_nativeaddress => nios2_clock_3_in_nativeaddress,
      nios2_clock_3_in_read => nios2_clock_3_in_read,
      nios2_clock_3_in_readdata_from_sa => nios2_clock_3_in_readdata_from_sa,
      nios2_clock_3_in_reset_n => nios2_clock_3_in_reset_n,
      nios2_clock_3_in_waitrequest_from_sa => nios2_clock_3_in_waitrequest_from_sa,
      nios2_clock_3_in_write => nios2_clock_3_in_write,
      nios2_clock_3_in_writedata => nios2_clock_3_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_3_in_endofpacket => nios2_clock_3_in_endofpacket,
      nios2_clock_3_in_readdata => nios2_clock_3_in_readdata,
      nios2_clock_3_in_waitrequest => nios2_clock_3_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_3_out, which is an e_instance
  the_nios2_clock_3_out : nios2_clock_3_out_arbitrator
    port map(
      nios2_clock_3_out_address_to_slave => nios2_clock_3_out_address_to_slave,
      nios2_clock_3_out_readdata => nios2_clock_3_out_readdata,
      nios2_clock_3_out_reset_n => nios2_clock_3_out_reset_n,
      nios2_clock_3_out_waitrequest => nios2_clock_3_out_waitrequest,
      clk => clk_0,
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      nios2_clock_3_out_address => nios2_clock_3_out_address,
      nios2_clock_3_out_byteenable => nios2_clock_3_out_byteenable,
      nios2_clock_3_out_granted_sys_clk_timer_s1 => nios2_clock_3_out_granted_sys_clk_timer_s1,
      nios2_clock_3_out_qualified_request_sys_clk_timer_s1 => nios2_clock_3_out_qualified_request_sys_clk_timer_s1,
      nios2_clock_3_out_read => nios2_clock_3_out_read,
      nios2_clock_3_out_read_data_valid_sys_clk_timer_s1 => nios2_clock_3_out_read_data_valid_sys_clk_timer_s1,
      nios2_clock_3_out_requests_sys_clk_timer_s1 => nios2_clock_3_out_requests_sys_clk_timer_s1,
      nios2_clock_3_out_write => nios2_clock_3_out_write,
      nios2_clock_3_out_writedata => nios2_clock_3_out_writedata,
      reset_n => clk_0_reset_n,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa
    );


  --the_nios2_clock_3, which is an e_ptf_instance
  the_nios2_clock_3 : nios2_clock_3
    port map(
      master_address => nios2_clock_3_out_address,
      master_byteenable => nios2_clock_3_out_byteenable,
      master_nativeaddress => nios2_clock_3_out_nativeaddress,
      master_read => nios2_clock_3_out_read,
      master_write => nios2_clock_3_out_write,
      master_writedata => nios2_clock_3_out_writedata,
      slave_endofpacket => nios2_clock_3_in_endofpacket,
      slave_readdata => nios2_clock_3_in_readdata,
      slave_waitrequest => nios2_clock_3_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_3_out_endofpacket,
      master_readdata => nios2_clock_3_out_readdata,
      master_reset_n => nios2_clock_3_out_reset_n,
      master_waitrequest => nios2_clock_3_out_waitrequest,
      slave_address => nios2_clock_3_in_address,
      slave_byteenable => nios2_clock_3_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_3_in_nativeaddress,
      slave_read => nios2_clock_3_in_read,
      slave_reset_n => nios2_clock_3_in_reset_n,
      slave_write => nios2_clock_3_in_write,
      slave_writedata => nios2_clock_3_in_writedata
    );


  --the_nios2_clock_4_in, which is an e_instance
  the_nios2_clock_4_in : nios2_clock_4_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_4_in => cpu_0_data_master_granted_nios2_clock_4_in,
      cpu_0_data_master_qualified_request_nios2_clock_4_in => cpu_0_data_master_qualified_request_nios2_clock_4_in,
      cpu_0_data_master_read_data_valid_nios2_clock_4_in => cpu_0_data_master_read_data_valid_nios2_clock_4_in,
      cpu_0_data_master_requests_nios2_clock_4_in => cpu_0_data_master_requests_nios2_clock_4_in,
      d1_nios2_clock_4_in_end_xfer => d1_nios2_clock_4_in_end_xfer,
      nios2_clock_4_in_address => nios2_clock_4_in_address,
      nios2_clock_4_in_byteenable => nios2_clock_4_in_byteenable,
      nios2_clock_4_in_endofpacket_from_sa => nios2_clock_4_in_endofpacket_from_sa,
      nios2_clock_4_in_nativeaddress => nios2_clock_4_in_nativeaddress,
      nios2_clock_4_in_read => nios2_clock_4_in_read,
      nios2_clock_4_in_readdata_from_sa => nios2_clock_4_in_readdata_from_sa,
      nios2_clock_4_in_reset_n => nios2_clock_4_in_reset_n,
      nios2_clock_4_in_waitrequest_from_sa => nios2_clock_4_in_waitrequest_from_sa,
      nios2_clock_4_in_write => nios2_clock_4_in_write,
      nios2_clock_4_in_writedata => nios2_clock_4_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_4_in_endofpacket => nios2_clock_4_in_endofpacket,
      nios2_clock_4_in_readdata => nios2_clock_4_in_readdata,
      nios2_clock_4_in_waitrequest => nios2_clock_4_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_4_out, which is an e_instance
  the_nios2_clock_4_out : nios2_clock_4_out_arbitrator
    port map(
      nios2_clock_4_out_address_to_slave => nios2_clock_4_out_address_to_slave,
      nios2_clock_4_out_readdata => nios2_clock_4_out_readdata,
      nios2_clock_4_out_reset_n => nios2_clock_4_out_reset_n,
      nios2_clock_4_out_waitrequest => nios2_clock_4_out_waitrequest,
      clk => clk_0,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      nios2_clock_4_out_address => nios2_clock_4_out_address,
      nios2_clock_4_out_byteenable => nios2_clock_4_out_byteenable,
      nios2_clock_4_out_granted_sysid_control_slave => nios2_clock_4_out_granted_sysid_control_slave,
      nios2_clock_4_out_qualified_request_sysid_control_slave => nios2_clock_4_out_qualified_request_sysid_control_slave,
      nios2_clock_4_out_read => nios2_clock_4_out_read,
      nios2_clock_4_out_read_data_valid_sysid_control_slave => nios2_clock_4_out_read_data_valid_sysid_control_slave,
      nios2_clock_4_out_requests_sysid_control_slave => nios2_clock_4_out_requests_sysid_control_slave,
      nios2_clock_4_out_write => nios2_clock_4_out_write,
      nios2_clock_4_out_writedata => nios2_clock_4_out_writedata,
      reset_n => clk_0_reset_n,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa
    );


  --the_nios2_clock_4, which is an e_ptf_instance
  the_nios2_clock_4 : nios2_clock_4
    port map(
      master_address => nios2_clock_4_out_address,
      master_byteenable => nios2_clock_4_out_byteenable,
      master_nativeaddress => nios2_clock_4_out_nativeaddress,
      master_read => nios2_clock_4_out_read,
      master_write => nios2_clock_4_out_write,
      master_writedata => nios2_clock_4_out_writedata,
      slave_endofpacket => nios2_clock_4_in_endofpacket,
      slave_readdata => nios2_clock_4_in_readdata,
      slave_waitrequest => nios2_clock_4_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_4_out_endofpacket,
      master_readdata => nios2_clock_4_out_readdata,
      master_reset_n => nios2_clock_4_out_reset_n,
      master_waitrequest => nios2_clock_4_out_waitrequest,
      slave_address => nios2_clock_4_in_address,
      slave_byteenable => nios2_clock_4_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_4_in_nativeaddress,
      slave_read => nios2_clock_4_in_read,
      slave_reset_n => nios2_clock_4_in_reset_n,
      slave_write => nios2_clock_4_in_write,
      slave_writedata => nios2_clock_4_in_writedata
    );


  --the_nios2_clock_5_in, which is an e_instance
  the_nios2_clock_5_in : nios2_clock_5_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_5_in => cpu_0_data_master_granted_nios2_clock_5_in,
      cpu_0_data_master_qualified_request_nios2_clock_5_in => cpu_0_data_master_qualified_request_nios2_clock_5_in,
      cpu_0_data_master_read_data_valid_nios2_clock_5_in => cpu_0_data_master_read_data_valid_nios2_clock_5_in,
      cpu_0_data_master_requests_nios2_clock_5_in => cpu_0_data_master_requests_nios2_clock_5_in,
      d1_nios2_clock_5_in_end_xfer => d1_nios2_clock_5_in_end_xfer,
      nios2_clock_5_in_address => nios2_clock_5_in_address,
      nios2_clock_5_in_byteenable => nios2_clock_5_in_byteenable,
      nios2_clock_5_in_endofpacket_from_sa => nios2_clock_5_in_endofpacket_from_sa,
      nios2_clock_5_in_nativeaddress => nios2_clock_5_in_nativeaddress,
      nios2_clock_5_in_read => nios2_clock_5_in_read,
      nios2_clock_5_in_readdata_from_sa => nios2_clock_5_in_readdata_from_sa,
      nios2_clock_5_in_reset_n => nios2_clock_5_in_reset_n,
      nios2_clock_5_in_waitrequest_from_sa => nios2_clock_5_in_waitrequest_from_sa,
      nios2_clock_5_in_write => nios2_clock_5_in_write,
      nios2_clock_5_in_writedata => nios2_clock_5_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_5_in_endofpacket => nios2_clock_5_in_endofpacket,
      nios2_clock_5_in_readdata => nios2_clock_5_in_readdata,
      nios2_clock_5_in_waitrequest => nios2_clock_5_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_5_out, which is an e_instance
  the_nios2_clock_5_out : nios2_clock_5_out_arbitrator
    port map(
      nios2_clock_5_out_address_to_slave => nios2_clock_5_out_address_to_slave,
      nios2_clock_5_out_readdata => nios2_clock_5_out_readdata,
      nios2_clock_5_out_reset_n => nios2_clock_5_out_reset_n,
      nios2_clock_5_out_waitrequest => nios2_clock_5_out_waitrequest,
      altpll_0_pll_slave_readdata_from_sa => altpll_0_pll_slave_readdata_from_sa,
      clk => clk_0,
      d1_altpll_0_pll_slave_end_xfer => d1_altpll_0_pll_slave_end_xfer,
      nios2_clock_5_out_address => nios2_clock_5_out_address,
      nios2_clock_5_out_byteenable => nios2_clock_5_out_byteenable,
      nios2_clock_5_out_granted_altpll_0_pll_slave => nios2_clock_5_out_granted_altpll_0_pll_slave,
      nios2_clock_5_out_qualified_request_altpll_0_pll_slave => nios2_clock_5_out_qualified_request_altpll_0_pll_slave,
      nios2_clock_5_out_read => nios2_clock_5_out_read,
      nios2_clock_5_out_read_data_valid_altpll_0_pll_slave => nios2_clock_5_out_read_data_valid_altpll_0_pll_slave,
      nios2_clock_5_out_requests_altpll_0_pll_slave => nios2_clock_5_out_requests_altpll_0_pll_slave,
      nios2_clock_5_out_write => nios2_clock_5_out_write,
      nios2_clock_5_out_writedata => nios2_clock_5_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_nios2_clock_5, which is an e_ptf_instance
  the_nios2_clock_5 : nios2_clock_5
    port map(
      master_address => nios2_clock_5_out_address,
      master_byteenable => nios2_clock_5_out_byteenable,
      master_nativeaddress => nios2_clock_5_out_nativeaddress,
      master_read => nios2_clock_5_out_read,
      master_write => nios2_clock_5_out_write,
      master_writedata => nios2_clock_5_out_writedata,
      slave_endofpacket => nios2_clock_5_in_endofpacket,
      slave_readdata => nios2_clock_5_in_readdata,
      slave_waitrequest => nios2_clock_5_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => nios2_clock_5_out_endofpacket,
      master_readdata => nios2_clock_5_out_readdata,
      master_reset_n => nios2_clock_5_out_reset_n,
      master_waitrequest => nios2_clock_5_out_waitrequest,
      slave_address => nios2_clock_5_in_address,
      slave_byteenable => nios2_clock_5_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_5_in_nativeaddress,
      slave_read => nios2_clock_5_in_read,
      slave_reset_n => nios2_clock_5_in_reset_n,
      slave_write => nios2_clock_5_in_write,
      slave_writedata => nios2_clock_5_in_writedata
    );


  --the_nios2_clock_6_in, which is an e_instance
  the_nios2_clock_6_in : nios2_clock_6_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_6_in => cpu_0_data_master_granted_nios2_clock_6_in,
      cpu_0_data_master_qualified_request_nios2_clock_6_in => cpu_0_data_master_qualified_request_nios2_clock_6_in,
      cpu_0_data_master_read_data_valid_nios2_clock_6_in => cpu_0_data_master_read_data_valid_nios2_clock_6_in,
      cpu_0_data_master_requests_nios2_clock_6_in => cpu_0_data_master_requests_nios2_clock_6_in,
      d1_nios2_clock_6_in_end_xfer => d1_nios2_clock_6_in_end_xfer,
      nios2_clock_6_in_address => nios2_clock_6_in_address,
      nios2_clock_6_in_byteenable => nios2_clock_6_in_byteenable,
      nios2_clock_6_in_endofpacket_from_sa => nios2_clock_6_in_endofpacket_from_sa,
      nios2_clock_6_in_nativeaddress => nios2_clock_6_in_nativeaddress,
      nios2_clock_6_in_read => nios2_clock_6_in_read,
      nios2_clock_6_in_readdata_from_sa => nios2_clock_6_in_readdata_from_sa,
      nios2_clock_6_in_reset_n => nios2_clock_6_in_reset_n,
      nios2_clock_6_in_waitrequest_from_sa => nios2_clock_6_in_waitrequest_from_sa,
      nios2_clock_6_in_write => nios2_clock_6_in_write,
      nios2_clock_6_in_writedata => nios2_clock_6_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_6_in_endofpacket => nios2_clock_6_in_endofpacket,
      nios2_clock_6_in_readdata => nios2_clock_6_in_readdata,
      nios2_clock_6_in_waitrequest => nios2_clock_6_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_6_out, which is an e_instance
  the_nios2_clock_6_out : nios2_clock_6_out_arbitrator
    port map(
      nios2_clock_6_out_address_to_slave => nios2_clock_6_out_address_to_slave,
      nios2_clock_6_out_readdata => nios2_clock_6_out_readdata,
      nios2_clock_6_out_reset_n => nios2_clock_6_out_reset_n,
      nios2_clock_6_out_waitrequest => nios2_clock_6_out_waitrequest,
      clk => internal_altpll_0_c0,
      d1_gen_code_value_pio_0_s1_end_xfer => d1_gen_code_value_pio_0_s1_end_xfer,
      gen_code_value_pio_0_s1_readdata_from_sa => gen_code_value_pio_0_s1_readdata_from_sa,
      nios2_clock_6_out_address => nios2_clock_6_out_address,
      nios2_clock_6_out_byteenable => nios2_clock_6_out_byteenable,
      nios2_clock_6_out_granted_gen_code_value_pio_0_s1 => nios2_clock_6_out_granted_gen_code_value_pio_0_s1,
      nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1 => nios2_clock_6_out_qualified_request_gen_code_value_pio_0_s1,
      nios2_clock_6_out_read => nios2_clock_6_out_read,
      nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1 => nios2_clock_6_out_read_data_valid_gen_code_value_pio_0_s1,
      nios2_clock_6_out_requests_gen_code_value_pio_0_s1 => nios2_clock_6_out_requests_gen_code_value_pio_0_s1,
      nios2_clock_6_out_write => nios2_clock_6_out_write,
      nios2_clock_6_out_writedata => nios2_clock_6_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_nios2_clock_6, which is an e_ptf_instance
  the_nios2_clock_6 : nios2_clock_6
    port map(
      master_address => nios2_clock_6_out_address,
      master_byteenable => nios2_clock_6_out_byteenable,
      master_nativeaddress => nios2_clock_6_out_nativeaddress,
      master_read => nios2_clock_6_out_read,
      master_write => nios2_clock_6_out_write,
      master_writedata => nios2_clock_6_out_writedata,
      slave_endofpacket => nios2_clock_6_in_endofpacket,
      slave_readdata => nios2_clock_6_in_readdata,
      slave_waitrequest => nios2_clock_6_in_waitrequest,
      master_clk => internal_altpll_0_c0,
      master_endofpacket => nios2_clock_6_out_endofpacket,
      master_readdata => nios2_clock_6_out_readdata,
      master_reset_n => nios2_clock_6_out_reset_n,
      master_waitrequest => nios2_clock_6_out_waitrequest,
      slave_address => nios2_clock_6_in_address,
      slave_byteenable => nios2_clock_6_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_6_in_nativeaddress,
      slave_read => nios2_clock_6_in_read,
      slave_reset_n => nios2_clock_6_in_reset_n,
      slave_write => nios2_clock_6_in_write,
      slave_writedata => nios2_clock_6_in_writedata
    );


  --the_nios2_clock_7_in, which is an e_instance
  the_nios2_clock_7_in : nios2_clock_7_in_arbitrator
    port map(
      cpu_0_data_master_granted_nios2_clock_7_in => cpu_0_data_master_granted_nios2_clock_7_in,
      cpu_0_data_master_qualified_request_nios2_clock_7_in => cpu_0_data_master_qualified_request_nios2_clock_7_in,
      cpu_0_data_master_read_data_valid_nios2_clock_7_in => cpu_0_data_master_read_data_valid_nios2_clock_7_in,
      cpu_0_data_master_requests_nios2_clock_7_in => cpu_0_data_master_requests_nios2_clock_7_in,
      d1_nios2_clock_7_in_end_xfer => d1_nios2_clock_7_in_end_xfer,
      nios2_clock_7_in_address => nios2_clock_7_in_address,
      nios2_clock_7_in_byteenable => nios2_clock_7_in_byteenable,
      nios2_clock_7_in_endofpacket_from_sa => nios2_clock_7_in_endofpacket_from_sa,
      nios2_clock_7_in_nativeaddress => nios2_clock_7_in_nativeaddress,
      nios2_clock_7_in_read => nios2_clock_7_in_read,
      nios2_clock_7_in_readdata_from_sa => nios2_clock_7_in_readdata_from_sa,
      nios2_clock_7_in_reset_n => nios2_clock_7_in_reset_n,
      nios2_clock_7_in_waitrequest_from_sa => nios2_clock_7_in_waitrequest_from_sa,
      nios2_clock_7_in_write => nios2_clock_7_in_write,
      nios2_clock_7_in_writedata => nios2_clock_7_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      nios2_clock_7_in_endofpacket => nios2_clock_7_in_endofpacket,
      nios2_clock_7_in_readdata => nios2_clock_7_in_readdata,
      nios2_clock_7_in_waitrequest => nios2_clock_7_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_7_out, which is an e_instance
  the_nios2_clock_7_out : nios2_clock_7_out_arbitrator
    port map(
      nios2_clock_7_out_address_to_slave => nios2_clock_7_out_address_to_slave,
      nios2_clock_7_out_readdata => nios2_clock_7_out_readdata,
      nios2_clock_7_out_reset_n => nios2_clock_7_out_reset_n,
      nios2_clock_7_out_waitrequest => nios2_clock_7_out_waitrequest,
      clk => internal_altpll_0_c0,
      d1_gen_code_value_pio_1_s1_end_xfer => d1_gen_code_value_pio_1_s1_end_xfer,
      gen_code_value_pio_1_s1_readdata_from_sa => gen_code_value_pio_1_s1_readdata_from_sa,
      nios2_clock_7_out_address => nios2_clock_7_out_address,
      nios2_clock_7_out_byteenable => nios2_clock_7_out_byteenable,
      nios2_clock_7_out_granted_gen_code_value_pio_1_s1 => nios2_clock_7_out_granted_gen_code_value_pio_1_s1,
      nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1 => nios2_clock_7_out_qualified_request_gen_code_value_pio_1_s1,
      nios2_clock_7_out_read => nios2_clock_7_out_read,
      nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1 => nios2_clock_7_out_read_data_valid_gen_code_value_pio_1_s1,
      nios2_clock_7_out_requests_gen_code_value_pio_1_s1 => nios2_clock_7_out_requests_gen_code_value_pio_1_s1,
      nios2_clock_7_out_write => nios2_clock_7_out_write,
      nios2_clock_7_out_writedata => nios2_clock_7_out_writedata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_nios2_clock_7, which is an e_ptf_instance
  the_nios2_clock_7 : nios2_clock_7
    port map(
      master_address => nios2_clock_7_out_address,
      master_byteenable => nios2_clock_7_out_byteenable,
      master_nativeaddress => nios2_clock_7_out_nativeaddress,
      master_read => nios2_clock_7_out_read,
      master_write => nios2_clock_7_out_write,
      master_writedata => nios2_clock_7_out_writedata,
      slave_endofpacket => nios2_clock_7_in_endofpacket,
      slave_readdata => nios2_clock_7_in_readdata,
      slave_waitrequest => nios2_clock_7_in_waitrequest,
      master_clk => internal_altpll_0_c0,
      master_endofpacket => nios2_clock_7_out_endofpacket,
      master_readdata => nios2_clock_7_out_readdata,
      master_reset_n => nios2_clock_7_out_reset_n,
      master_waitrequest => nios2_clock_7_out_waitrequest,
      slave_address => nios2_clock_7_in_address,
      slave_byteenable => nios2_clock_7_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_7_in_nativeaddress,
      slave_read => nios2_clock_7_in_read,
      slave_reset_n => nios2_clock_7_in_reset_n,
      slave_write => nios2_clock_7_in_write,
      slave_writedata => nios2_clock_7_in_writedata
    );


  --the_nios2_clock_8_in, which is an e_instance
  the_nios2_clock_8_in : nios2_clock_8_in_arbitrator
    port map(
      cpu_0_instruction_master_granted_nios2_clock_8_in => cpu_0_instruction_master_granted_nios2_clock_8_in,
      cpu_0_instruction_master_qualified_request_nios2_clock_8_in => cpu_0_instruction_master_qualified_request_nios2_clock_8_in,
      cpu_0_instruction_master_read_data_valid_nios2_clock_8_in => cpu_0_instruction_master_read_data_valid_nios2_clock_8_in,
      cpu_0_instruction_master_requests_nios2_clock_8_in => cpu_0_instruction_master_requests_nios2_clock_8_in,
      d1_nios2_clock_8_in_end_xfer => d1_nios2_clock_8_in_end_xfer,
      nios2_clock_8_in_address => nios2_clock_8_in_address,
      nios2_clock_8_in_byteenable => nios2_clock_8_in_byteenable,
      nios2_clock_8_in_endofpacket_from_sa => nios2_clock_8_in_endofpacket_from_sa,
      nios2_clock_8_in_nativeaddress => nios2_clock_8_in_nativeaddress,
      nios2_clock_8_in_read => nios2_clock_8_in_read,
      nios2_clock_8_in_readdata_from_sa => nios2_clock_8_in_readdata_from_sa,
      nios2_clock_8_in_reset_n => nios2_clock_8_in_reset_n,
      nios2_clock_8_in_waitrequest_from_sa => nios2_clock_8_in_waitrequest_from_sa,
      nios2_clock_8_in_write => nios2_clock_8_in_write,
      clk => processor_clk,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_dbs_address => cpu_0_instruction_master_dbs_address,
      cpu_0_instruction_master_latency_counter => cpu_0_instruction_master_latency_counter,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      nios2_clock_8_in_endofpacket => nios2_clock_8_in_endofpacket,
      nios2_clock_8_in_readdata => nios2_clock_8_in_readdata,
      nios2_clock_8_in_waitrequest => nios2_clock_8_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_8_out, which is an e_instance
  the_nios2_clock_8_out : nios2_clock_8_out_arbitrator
    port map(
      nios2_clock_8_out_address_to_slave => nios2_clock_8_out_address_to_slave,
      nios2_clock_8_out_readdata => nios2_clock_8_out_readdata,
      nios2_clock_8_out_reset_n => nios2_clock_8_out_reset_n,
      nios2_clock_8_out_waitrequest => nios2_clock_8_out_waitrequest,
      clk => internal_altpll_0_c1_out,
      d1_sdram_0_s1_end_xfer => d1_sdram_0_s1_end_xfer,
      nios2_clock_8_out_address => nios2_clock_8_out_address,
      nios2_clock_8_out_byteenable => nios2_clock_8_out_byteenable,
      nios2_clock_8_out_granted_sdram_0_s1 => nios2_clock_8_out_granted_sdram_0_s1,
      nios2_clock_8_out_qualified_request_sdram_0_s1 => nios2_clock_8_out_qualified_request_sdram_0_s1,
      nios2_clock_8_out_read => nios2_clock_8_out_read,
      nios2_clock_8_out_read_data_valid_sdram_0_s1 => nios2_clock_8_out_read_data_valid_sdram_0_s1,
      nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register => nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register,
      nios2_clock_8_out_requests_sdram_0_s1 => nios2_clock_8_out_requests_sdram_0_s1,
      nios2_clock_8_out_write => nios2_clock_8_out_write,
      nios2_clock_8_out_writedata => nios2_clock_8_out_writedata,
      reset_n => altpll_0_c1_out_reset_n,
      sdram_0_s1_readdata_from_sa => sdram_0_s1_readdata_from_sa,
      sdram_0_s1_waitrequest_from_sa => sdram_0_s1_waitrequest_from_sa
    );


  --the_nios2_clock_8, which is an e_ptf_instance
  the_nios2_clock_8 : nios2_clock_8
    port map(
      master_address => nios2_clock_8_out_address,
      master_byteenable => nios2_clock_8_out_byteenable,
      master_nativeaddress => nios2_clock_8_out_nativeaddress,
      master_read => nios2_clock_8_out_read,
      master_write => nios2_clock_8_out_write,
      master_writedata => nios2_clock_8_out_writedata,
      slave_endofpacket => nios2_clock_8_in_endofpacket,
      slave_readdata => nios2_clock_8_in_readdata,
      slave_waitrequest => nios2_clock_8_in_waitrequest,
      master_clk => internal_altpll_0_c1_out,
      master_endofpacket => nios2_clock_8_out_endofpacket,
      master_readdata => nios2_clock_8_out_readdata,
      master_reset_n => nios2_clock_8_out_reset_n,
      master_waitrequest => nios2_clock_8_out_waitrequest,
      slave_address => nios2_clock_8_in_address,
      slave_byteenable => nios2_clock_8_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_8_in_nativeaddress,
      slave_read => nios2_clock_8_in_read,
      slave_reset_n => nios2_clock_8_in_reset_n,
      slave_write => nios2_clock_8_in_write,
      slave_writedata => nios2_clock_8_in_writedata
    );


  --the_nios2_clock_9_in, which is an e_instance
  the_nios2_clock_9_in : nios2_clock_9_in_arbitrator
    port map(
      cpu_0_data_master_byteenable_nios2_clock_9_in => cpu_0_data_master_byteenable_nios2_clock_9_in,
      cpu_0_data_master_granted_nios2_clock_9_in => cpu_0_data_master_granted_nios2_clock_9_in,
      cpu_0_data_master_qualified_request_nios2_clock_9_in => cpu_0_data_master_qualified_request_nios2_clock_9_in,
      cpu_0_data_master_read_data_valid_nios2_clock_9_in => cpu_0_data_master_read_data_valid_nios2_clock_9_in,
      cpu_0_data_master_requests_nios2_clock_9_in => cpu_0_data_master_requests_nios2_clock_9_in,
      d1_nios2_clock_9_in_end_xfer => d1_nios2_clock_9_in_end_xfer,
      nios2_clock_9_in_address => nios2_clock_9_in_address,
      nios2_clock_9_in_byteenable => nios2_clock_9_in_byteenable,
      nios2_clock_9_in_endofpacket_from_sa => nios2_clock_9_in_endofpacket_from_sa,
      nios2_clock_9_in_nativeaddress => nios2_clock_9_in_nativeaddress,
      nios2_clock_9_in_read => nios2_clock_9_in_read,
      nios2_clock_9_in_readdata_from_sa => nios2_clock_9_in_readdata_from_sa,
      nios2_clock_9_in_reset_n => nios2_clock_9_in_reset_n,
      nios2_clock_9_in_waitrequest_from_sa => nios2_clock_9_in_waitrequest_from_sa,
      nios2_clock_9_in_write => nios2_clock_9_in_write,
      nios2_clock_9_in_writedata => nios2_clock_9_in_writedata,
      clk => processor_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_dbs_address => cpu_0_data_master_dbs_address,
      cpu_0_data_master_dbs_write_16 => cpu_0_data_master_dbs_write_16,
      cpu_0_data_master_latency_counter => cpu_0_data_master_latency_counter,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_write => cpu_0_data_master_write,
      nios2_clock_9_in_endofpacket => nios2_clock_9_in_endofpacket,
      nios2_clock_9_in_readdata => nios2_clock_9_in_readdata,
      nios2_clock_9_in_waitrequest => nios2_clock_9_in_waitrequest,
      reset_n => processor_clk_reset_n
    );


  --the_nios2_clock_9_out, which is an e_instance
  the_nios2_clock_9_out : nios2_clock_9_out_arbitrator
    port map(
      nios2_clock_9_out_address_to_slave => nios2_clock_9_out_address_to_slave,
      nios2_clock_9_out_readdata => nios2_clock_9_out_readdata,
      nios2_clock_9_out_reset_n => nios2_clock_9_out_reset_n,
      nios2_clock_9_out_waitrequest => nios2_clock_9_out_waitrequest,
      clk => internal_altpll_0_c1_out,
      d1_sdram_0_s1_end_xfer => d1_sdram_0_s1_end_xfer,
      nios2_clock_9_out_address => nios2_clock_9_out_address,
      nios2_clock_9_out_byteenable => nios2_clock_9_out_byteenable,
      nios2_clock_9_out_granted_sdram_0_s1 => nios2_clock_9_out_granted_sdram_0_s1,
      nios2_clock_9_out_qualified_request_sdram_0_s1 => nios2_clock_9_out_qualified_request_sdram_0_s1,
      nios2_clock_9_out_read => nios2_clock_9_out_read,
      nios2_clock_9_out_read_data_valid_sdram_0_s1 => nios2_clock_9_out_read_data_valid_sdram_0_s1,
      nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register => nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register,
      nios2_clock_9_out_requests_sdram_0_s1 => nios2_clock_9_out_requests_sdram_0_s1,
      nios2_clock_9_out_write => nios2_clock_9_out_write,
      nios2_clock_9_out_writedata => nios2_clock_9_out_writedata,
      reset_n => altpll_0_c1_out_reset_n,
      sdram_0_s1_readdata_from_sa => sdram_0_s1_readdata_from_sa,
      sdram_0_s1_waitrequest_from_sa => sdram_0_s1_waitrequest_from_sa
    );


  --the_nios2_clock_9, which is an e_ptf_instance
  the_nios2_clock_9 : nios2_clock_9
    port map(
      master_address => nios2_clock_9_out_address,
      master_byteenable => nios2_clock_9_out_byteenable,
      master_nativeaddress => nios2_clock_9_out_nativeaddress,
      master_read => nios2_clock_9_out_read,
      master_write => nios2_clock_9_out_write,
      master_writedata => nios2_clock_9_out_writedata,
      slave_endofpacket => nios2_clock_9_in_endofpacket,
      slave_readdata => nios2_clock_9_in_readdata,
      slave_waitrequest => nios2_clock_9_in_waitrequest,
      master_clk => internal_altpll_0_c1_out,
      master_endofpacket => nios2_clock_9_out_endofpacket,
      master_readdata => nios2_clock_9_out_readdata,
      master_reset_n => nios2_clock_9_out_reset_n,
      master_waitrequest => nios2_clock_9_out_waitrequest,
      slave_address => nios2_clock_9_in_address,
      slave_byteenable => nios2_clock_9_in_byteenable,
      slave_clk => processor_clk,
      slave_nativeaddress => nios2_clock_9_in_nativeaddress,
      slave_read => nios2_clock_9_in_read,
      slave_reset_n => nios2_clock_9_in_reset_n,
      slave_write => nios2_clock_9_in_write,
      slave_writedata => nios2_clock_9_in_writedata
    );


  --the_onchip_mem_s1, which is an e_instance
  the_onchip_mem_s1 : onchip_mem_s1_arbitrator
    port map(
      d1_onchip_mem_s1_end_xfer => d1_onchip_mem_s1_end_xfer,
      nios2_clock_0_out_granted_onchip_mem_s1 => nios2_clock_0_out_granted_onchip_mem_s1,
      nios2_clock_0_out_qualified_request_onchip_mem_s1 => nios2_clock_0_out_qualified_request_onchip_mem_s1,
      nios2_clock_0_out_read_data_valid_onchip_mem_s1 => nios2_clock_0_out_read_data_valid_onchip_mem_s1,
      nios2_clock_0_out_requests_onchip_mem_s1 => nios2_clock_0_out_requests_onchip_mem_s1,
      nios2_clock_1_out_granted_onchip_mem_s1 => nios2_clock_1_out_granted_onchip_mem_s1,
      nios2_clock_1_out_qualified_request_onchip_mem_s1 => nios2_clock_1_out_qualified_request_onchip_mem_s1,
      nios2_clock_1_out_read_data_valid_onchip_mem_s1 => nios2_clock_1_out_read_data_valid_onchip_mem_s1,
      nios2_clock_1_out_requests_onchip_mem_s1 => nios2_clock_1_out_requests_onchip_mem_s1,
      onchip_mem_s1_address => onchip_mem_s1_address,
      onchip_mem_s1_byteenable => onchip_mem_s1_byteenable,
      onchip_mem_s1_chipselect => onchip_mem_s1_chipselect,
      onchip_mem_s1_clken => onchip_mem_s1_clken,
      onchip_mem_s1_readdata_from_sa => onchip_mem_s1_readdata_from_sa,
      onchip_mem_s1_reset => onchip_mem_s1_reset,
      onchip_mem_s1_write => onchip_mem_s1_write,
      onchip_mem_s1_writedata => onchip_mem_s1_writedata,
      clk => internal_altpll_0_c0,
      nios2_clock_0_out_address_to_slave => nios2_clock_0_out_address_to_slave,
      nios2_clock_0_out_byteenable => nios2_clock_0_out_byteenable,
      nios2_clock_0_out_read => nios2_clock_0_out_read,
      nios2_clock_0_out_write => nios2_clock_0_out_write,
      nios2_clock_0_out_writedata => nios2_clock_0_out_writedata,
      nios2_clock_1_out_address_to_slave => nios2_clock_1_out_address_to_slave,
      nios2_clock_1_out_byteenable => nios2_clock_1_out_byteenable,
      nios2_clock_1_out_read => nios2_clock_1_out_read,
      nios2_clock_1_out_write => nios2_clock_1_out_write,
      nios2_clock_1_out_writedata => nios2_clock_1_out_writedata,
      onchip_mem_s1_readdata => onchip_mem_s1_readdata,
      reset_n => altpll_0_c0_reset_n
    );


  --the_onchip_mem, which is an e_ptf_instance
  the_onchip_mem : onchip_mem
    port map(
      readdata => onchip_mem_s1_readdata,
      address => onchip_mem_s1_address,
      byteenable => onchip_mem_s1_byteenable,
      chipselect => onchip_mem_s1_chipselect,
      clk => internal_altpll_0_c0,
      clken => onchip_mem_s1_clken,
      reset => onchip_mem_s1_reset,
      write => onchip_mem_s1_write,
      writedata => onchip_mem_s1_writedata
    );


  --the_sample_and_hold_pio_s1, which is an e_instance
  the_sample_and_hold_pio_s1 : sample_and_hold_pio_s1_arbitrator
    port map(
      d1_sample_and_hold_pio_s1_end_xfer => d1_sample_and_hold_pio_s1_end_xfer,
      nios2_clock_17_out_granted_sample_and_hold_pio_s1 => nios2_clock_17_out_granted_sample_and_hold_pio_s1,
      nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1 => nios2_clock_17_out_qualified_request_sample_and_hold_pio_s1,
      nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1 => nios2_clock_17_out_read_data_valid_sample_and_hold_pio_s1,
      nios2_clock_17_out_requests_sample_and_hold_pio_s1 => nios2_clock_17_out_requests_sample_and_hold_pio_s1,
      sample_and_hold_pio_s1_address => sample_and_hold_pio_s1_address,
      sample_and_hold_pio_s1_chipselect => sample_and_hold_pio_s1_chipselect,
      sample_and_hold_pio_s1_readdata_from_sa => sample_and_hold_pio_s1_readdata_from_sa,
      sample_and_hold_pio_s1_reset_n => sample_and_hold_pio_s1_reset_n,
      sample_and_hold_pio_s1_write_n => sample_and_hold_pio_s1_write_n,
      sample_and_hold_pio_s1_writedata => sample_and_hold_pio_s1_writedata,
      clk => clk_0,
      nios2_clock_17_out_address_to_slave => nios2_clock_17_out_address_to_slave,
      nios2_clock_17_out_nativeaddress => nios2_clock_17_out_nativeaddress,
      nios2_clock_17_out_read => nios2_clock_17_out_read,
      nios2_clock_17_out_write => nios2_clock_17_out_write,
      nios2_clock_17_out_writedata => nios2_clock_17_out_writedata,
      reset_n => clk_0_reset_n,
      sample_and_hold_pio_s1_readdata => sample_and_hold_pio_s1_readdata
    );


  --the_sample_and_hold_pio, which is an e_ptf_instance
  the_sample_and_hold_pio : sample_and_hold_pio
    port map(
      out_port => internal_out_port_from_the_sample_and_hold_pio,
      readdata => sample_and_hold_pio_s1_readdata,
      address => sample_and_hold_pio_s1_address,
      chipselect => sample_and_hold_pio_s1_chipselect,
      clk => clk_0,
      reset_n => sample_and_hold_pio_s1_reset_n,
      write_n => sample_and_hold_pio_s1_write_n,
      writedata => sample_and_hold_pio_s1_writedata
    );


  --the_sdram_0_s1, which is an e_instance
  the_sdram_0_s1 : sdram_0_s1_arbitrator
    port map(
      d1_sdram_0_s1_end_xfer => d1_sdram_0_s1_end_xfer,
      nios2_clock_8_out_granted_sdram_0_s1 => nios2_clock_8_out_granted_sdram_0_s1,
      nios2_clock_8_out_qualified_request_sdram_0_s1 => nios2_clock_8_out_qualified_request_sdram_0_s1,
      nios2_clock_8_out_read_data_valid_sdram_0_s1 => nios2_clock_8_out_read_data_valid_sdram_0_s1,
      nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register => nios2_clock_8_out_read_data_valid_sdram_0_s1_shift_register,
      nios2_clock_8_out_requests_sdram_0_s1 => nios2_clock_8_out_requests_sdram_0_s1,
      nios2_clock_9_out_granted_sdram_0_s1 => nios2_clock_9_out_granted_sdram_0_s1,
      nios2_clock_9_out_qualified_request_sdram_0_s1 => nios2_clock_9_out_qualified_request_sdram_0_s1,
      nios2_clock_9_out_read_data_valid_sdram_0_s1 => nios2_clock_9_out_read_data_valid_sdram_0_s1,
      nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register => nios2_clock_9_out_read_data_valid_sdram_0_s1_shift_register,
      nios2_clock_9_out_requests_sdram_0_s1 => nios2_clock_9_out_requests_sdram_0_s1,
      sdram_0_s1_address => sdram_0_s1_address,
      sdram_0_s1_byteenable_n => sdram_0_s1_byteenable_n,
      sdram_0_s1_chipselect => sdram_0_s1_chipselect,
      sdram_0_s1_read_n => sdram_0_s1_read_n,
      sdram_0_s1_readdata_from_sa => sdram_0_s1_readdata_from_sa,
      sdram_0_s1_reset_n => sdram_0_s1_reset_n,
      sdram_0_s1_waitrequest_from_sa => sdram_0_s1_waitrequest_from_sa,
      sdram_0_s1_write_n => sdram_0_s1_write_n,
      sdram_0_s1_writedata => sdram_0_s1_writedata,
      clk => internal_altpll_0_c1_out,
      nios2_clock_8_out_address_to_slave => nios2_clock_8_out_address_to_slave,
      nios2_clock_8_out_byteenable => nios2_clock_8_out_byteenable,
      nios2_clock_8_out_read => nios2_clock_8_out_read,
      nios2_clock_8_out_write => nios2_clock_8_out_write,
      nios2_clock_8_out_writedata => nios2_clock_8_out_writedata,
      nios2_clock_9_out_address_to_slave => nios2_clock_9_out_address_to_slave,
      nios2_clock_9_out_byteenable => nios2_clock_9_out_byteenable,
      nios2_clock_9_out_read => nios2_clock_9_out_read,
      nios2_clock_9_out_write => nios2_clock_9_out_write,
      nios2_clock_9_out_writedata => nios2_clock_9_out_writedata,
      reset_n => altpll_0_c1_out_reset_n,
      sdram_0_s1_readdata => sdram_0_s1_readdata,
      sdram_0_s1_readdatavalid => sdram_0_s1_readdatavalid,
      sdram_0_s1_waitrequest => sdram_0_s1_waitrequest
    );


  --the_sdram_0, which is an e_ptf_instance
  the_sdram_0 : sdram_0
    port map(
      za_data => sdram_0_s1_readdata,
      za_valid => sdram_0_s1_readdatavalid,
      za_waitrequest => sdram_0_s1_waitrequest,
      zs_addr => internal_zs_addr_from_the_sdram_0,
      zs_ba => internal_zs_ba_from_the_sdram_0,
      zs_cas_n => internal_zs_cas_n_from_the_sdram_0,
      zs_cke => internal_zs_cke_from_the_sdram_0,
      zs_cs_n => internal_zs_cs_n_from_the_sdram_0,
      zs_dq => zs_dq_to_and_from_the_sdram_0,
      zs_dqm => internal_zs_dqm_from_the_sdram_0,
      zs_ras_n => internal_zs_ras_n_from_the_sdram_0,
      zs_we_n => internal_zs_we_n_from_the_sdram_0,
      az_addr => sdram_0_s1_address,
      az_be_n => sdram_0_s1_byteenable_n,
      az_cs => sdram_0_s1_chipselect,
      az_data => sdram_0_s1_writedata,
      az_rd_n => sdram_0_s1_read_n,
      az_wr_n => sdram_0_s1_write_n,
      clk => internal_altpll_0_c1_out,
      reset_n => sdram_0_s1_reset_n
    );


  --the_switch_pio_s1, which is an e_instance
  the_switch_pio_s1 : switch_pio_s1_arbitrator
    port map(
      d1_switch_pio_s1_end_xfer => d1_switch_pio_s1_end_xfer,
      nios2_clock_14_out_granted_switch_pio_s1 => nios2_clock_14_out_granted_switch_pio_s1,
      nios2_clock_14_out_qualified_request_switch_pio_s1 => nios2_clock_14_out_qualified_request_switch_pio_s1,
      nios2_clock_14_out_read_data_valid_switch_pio_s1 => nios2_clock_14_out_read_data_valid_switch_pio_s1,
      nios2_clock_14_out_requests_switch_pio_s1 => nios2_clock_14_out_requests_switch_pio_s1,
      switch_pio_s1_address => switch_pio_s1_address,
      switch_pio_s1_chipselect => switch_pio_s1_chipselect,
      switch_pio_s1_readdata_from_sa => switch_pio_s1_readdata_from_sa,
      switch_pio_s1_reset_n => switch_pio_s1_reset_n,
      switch_pio_s1_write_n => switch_pio_s1_write_n,
      switch_pio_s1_writedata => switch_pio_s1_writedata,
      clk => clk_0,
      nios2_clock_14_out_address_to_slave => nios2_clock_14_out_address_to_slave,
      nios2_clock_14_out_nativeaddress => nios2_clock_14_out_nativeaddress,
      nios2_clock_14_out_read => nios2_clock_14_out_read,
      nios2_clock_14_out_write => nios2_clock_14_out_write,
      nios2_clock_14_out_writedata => nios2_clock_14_out_writedata,
      reset_n => clk_0_reset_n,
      switch_pio_s1_readdata => switch_pio_s1_readdata
    );


  --the_switch_pio, which is an e_ptf_instance
  the_switch_pio : switch_pio
    port map(
      out_port => internal_out_port_from_the_switch_pio,
      readdata => switch_pio_s1_readdata,
      address => switch_pio_s1_address,
      chipselect => switch_pio_s1_chipselect,
      clk => clk_0,
      reset_n => switch_pio_s1_reset_n,
      write_n => switch_pio_s1_write_n,
      writedata => switch_pio_s1_writedata
    );


  --the_sys_clk_timer_s1, which is an e_instance
  the_sys_clk_timer_s1 : sys_clk_timer_s1_arbitrator
    port map(
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      nios2_clock_3_out_granted_sys_clk_timer_s1 => nios2_clock_3_out_granted_sys_clk_timer_s1,
      nios2_clock_3_out_qualified_request_sys_clk_timer_s1 => nios2_clock_3_out_qualified_request_sys_clk_timer_s1,
      nios2_clock_3_out_read_data_valid_sys_clk_timer_s1 => nios2_clock_3_out_read_data_valid_sys_clk_timer_s1,
      nios2_clock_3_out_requests_sys_clk_timer_s1 => nios2_clock_3_out_requests_sys_clk_timer_s1,
      sys_clk_timer_s1_address => sys_clk_timer_s1_address,
      sys_clk_timer_s1_chipselect => sys_clk_timer_s1_chipselect,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa,
      sys_clk_timer_s1_reset_n => sys_clk_timer_s1_reset_n,
      sys_clk_timer_s1_write_n => sys_clk_timer_s1_write_n,
      sys_clk_timer_s1_writedata => sys_clk_timer_s1_writedata,
      clk => clk_0,
      nios2_clock_3_out_address_to_slave => nios2_clock_3_out_address_to_slave,
      nios2_clock_3_out_nativeaddress => nios2_clock_3_out_nativeaddress,
      nios2_clock_3_out_read => nios2_clock_3_out_read,
      nios2_clock_3_out_write => nios2_clock_3_out_write,
      nios2_clock_3_out_writedata => nios2_clock_3_out_writedata,
      reset_n => clk_0_reset_n,
      sys_clk_timer_s1_irq => sys_clk_timer_s1_irq,
      sys_clk_timer_s1_readdata => sys_clk_timer_s1_readdata
    );


  --the_sys_clk_timer, which is an e_ptf_instance
  the_sys_clk_timer : sys_clk_timer
    port map(
      irq => sys_clk_timer_s1_irq,
      readdata => sys_clk_timer_s1_readdata,
      address => sys_clk_timer_s1_address,
      chipselect => sys_clk_timer_s1_chipselect,
      clk => clk_0,
      reset_n => sys_clk_timer_s1_reset_n,
      write_n => sys_clk_timer_s1_write_n,
      writedata => sys_clk_timer_s1_writedata
    );


  --the_sysid_control_slave, which is an e_instance
  the_sysid_control_slave : sysid_control_slave_arbitrator
    port map(
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      nios2_clock_4_out_granted_sysid_control_slave => nios2_clock_4_out_granted_sysid_control_slave,
      nios2_clock_4_out_qualified_request_sysid_control_slave => nios2_clock_4_out_qualified_request_sysid_control_slave,
      nios2_clock_4_out_read_data_valid_sysid_control_slave => nios2_clock_4_out_read_data_valid_sysid_control_slave,
      nios2_clock_4_out_requests_sysid_control_slave => nios2_clock_4_out_requests_sysid_control_slave,
      sysid_control_slave_address => sysid_control_slave_address,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      sysid_control_slave_reset_n => sysid_control_slave_reset_n,
      clk => clk_0,
      nios2_clock_4_out_address_to_slave => nios2_clock_4_out_address_to_slave,
      nios2_clock_4_out_nativeaddress => nios2_clock_4_out_nativeaddress,
      nios2_clock_4_out_read => nios2_clock_4_out_read,
      nios2_clock_4_out_write => nios2_clock_4_out_write,
      reset_n => clk_0_reset_n,
      sysid_control_slave_readdata => sysid_control_slave_readdata
    );


  --the_sysid, which is an e_ptf_instance
  the_sysid : sysid
    port map(
      readdata => sysid_control_slave_readdata,
      address => sysid_control_slave_address,
      clock => sysid_control_slave_clock,
      reset_n => sysid_control_slave_reset_n
    );


  --the_usb_code_pio_s1, which is an e_instance
  the_usb_code_pio_s1 : usb_code_pio_s1_arbitrator
    port map(
      d1_usb_code_pio_s1_end_xfer => d1_usb_code_pio_s1_end_xfer,
      nios2_clock_16_out_granted_usb_code_pio_s1 => nios2_clock_16_out_granted_usb_code_pio_s1,
      nios2_clock_16_out_qualified_request_usb_code_pio_s1 => nios2_clock_16_out_qualified_request_usb_code_pio_s1,
      nios2_clock_16_out_read_data_valid_usb_code_pio_s1 => nios2_clock_16_out_read_data_valid_usb_code_pio_s1,
      nios2_clock_16_out_requests_usb_code_pio_s1 => nios2_clock_16_out_requests_usb_code_pio_s1,
      usb_code_pio_s1_address => usb_code_pio_s1_address,
      usb_code_pio_s1_chipselect => usb_code_pio_s1_chipselect,
      usb_code_pio_s1_readdata_from_sa => usb_code_pio_s1_readdata_from_sa,
      usb_code_pio_s1_reset_n => usb_code_pio_s1_reset_n,
      usb_code_pio_s1_write_n => usb_code_pio_s1_write_n,
      usb_code_pio_s1_writedata => usb_code_pio_s1_writedata,
      clk => clk_0,
      nios2_clock_16_out_address_to_slave => nios2_clock_16_out_address_to_slave,
      nios2_clock_16_out_nativeaddress => nios2_clock_16_out_nativeaddress,
      nios2_clock_16_out_read => nios2_clock_16_out_read,
      nios2_clock_16_out_write => nios2_clock_16_out_write,
      nios2_clock_16_out_writedata => nios2_clock_16_out_writedata,
      reset_n => clk_0_reset_n,
      usb_code_pio_s1_readdata => usb_code_pio_s1_readdata
    );


  --the_usb_code_pio, which is an e_ptf_instance
  the_usb_code_pio : usb_code_pio
    port map(
      out_port => internal_out_port_from_the_usb_code_pio,
      readdata => usb_code_pio_s1_readdata,
      address => usb_code_pio_s1_address,
      chipselect => usb_code_pio_s1_chipselect,
      clk => clk_0,
      reset_n => usb_code_pio_s1_reset_n,
      write_n => usb_code_pio_s1_write_n,
      writedata => usb_code_pio_s1_writedata
    );


  --reset is asserted asynchronously and deasserted synchronously
  nios2_reset_clk_0_domain_synch : nios2_reset_clk_0_domain_synch_module
    port map(
      data_out => clk_0_reset_n,
      clk => clk_0,
      data_in => module_input6,
      reset_n => reset_n_sources
    );

  module_input6 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT ((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000"))));
  --reset is asserted asynchronously and deasserted synchronously
  nios2_reset_altpll_0_c0_domain_synch : nios2_reset_altpll_0_c0_domain_synch_module
    port map(
      data_out => altpll_0_c0_reset_n,
      clk => internal_altpll_0_c0,
      data_in => module_input7,
      reset_n => reset_n_sources
    );

  module_input7 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  nios2_reset_processor_clk_domain_synch : nios2_reset_processor_clk_domain_synch_module
    port map(
      data_out => processor_clk_reset_n,
      clk => processor_clk,
      data_in => module_input8,
      reset_n => reset_n_sources
    );

  module_input8 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  nios2_reset_altpll_0_c1_out_domain_synch : nios2_reset_altpll_0_c1_out_domain_synch_module
    port map(
      data_out => altpll_0_c1_out_reset_n,
      clk => internal_altpll_0_c1_out,
      data_in => module_input9,
      reset_n => reset_n_sources
    );

  module_input9 <= std_logic'('1');

  --nios2_clock_0_in_writedata of type writedata does not connect to anything so wire it to default (0)
  nios2_clock_0_in_writedata <= std_logic_vector'("00000000000000000000000000000000");
  --nios2_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_0_out_endofpacket <= std_logic'('0');
  --nios2_clock_10_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_10_out_endofpacket <= std_logic'('0');
  --nios2_clock_11_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_11_out_endofpacket <= std_logic'('0');
  --nios2_clock_12_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_12_out_endofpacket <= std_logic'('0');
  --nios2_clock_13_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_13_out_endofpacket <= std_logic'('0');
  --nios2_clock_14_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_14_out_endofpacket <= std_logic'('0');
  --nios2_clock_15_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_15_out_endofpacket <= std_logic'('0');
  --nios2_clock_16_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_16_out_endofpacket <= std_logic'('0');
  --nios2_clock_17_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_17_out_endofpacket <= std_logic'('0');
  --nios2_clock_18_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_18_out_endofpacket <= std_logic'('0');
  --nios2_clock_1_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_1_out_endofpacket <= std_logic'('0');
  --nios2_clock_2_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_2_out_endofpacket <= std_logic'('0');
  --nios2_clock_3_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_3_out_endofpacket <= std_logic'('0');
  --nios2_clock_4_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_4_out_endofpacket <= std_logic'('0');
  --nios2_clock_5_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_5_out_endofpacket <= std_logic'('0');
  --nios2_clock_6_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_6_out_endofpacket <= std_logic'('0');
  --nios2_clock_7_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_7_out_endofpacket <= std_logic'('0');
  --nios2_clock_8_in_writedata of type writedata does not connect to anything so wire it to default (0)
  nios2_clock_8_in_writedata <= std_logic_vector'("0000000000000000");
  --nios2_clock_8_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_8_out_endofpacket <= std_logic'('0');
  --nios2_clock_9_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  nios2_clock_9_out_endofpacket <= std_logic'('0');
  --sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  sysid_control_slave_clock <= std_logic'('0');
  --vhdl renameroo for output signals
  altpll_0_c0 <= internal_altpll_0_c0;
  --vhdl renameroo for output signals
  altpll_0_c1_out <= internal_altpll_0_c1_out;
  --vhdl renameroo for output signals
  locked_from_the_altpll_0 <= internal_locked_from_the_altpll_0;
  --vhdl renameroo for output signals
  out_port_from_the_cal_dac_code_pio <= internal_out_port_from_the_cal_dac_code_pio;
  --vhdl renameroo for output signals
  out_port_from_the_gen_code_strobe <= internal_out_port_from_the_gen_code_strobe;
  --vhdl renameroo for output signals
  out_port_from_the_gen_code_value_pio_0 <= internal_out_port_from_the_gen_code_value_pio_0;
  --vhdl renameroo for output signals
  out_port_from_the_gen_code_value_pio_1 <= internal_out_port_from_the_gen_code_value_pio_1;
  --vhdl renameroo for output signals
  out_port_from_the_latch_pio <= internal_out_port_from_the_latch_pio;
  --vhdl renameroo for output signals
  out_port_from_the_led_pio <= internal_out_port_from_the_led_pio;
  --vhdl renameroo for output signals
  out_port_from_the_sample_and_hold_pio <= internal_out_port_from_the_sample_and_hold_pio;
  --vhdl renameroo for output signals
  out_port_from_the_switch_pio <= internal_out_port_from_the_switch_pio;
  --vhdl renameroo for output signals
  out_port_from_the_usb_code_pio <= internal_out_port_from_the_usb_code_pio;
  --vhdl renameroo for output signals
  phasedone_from_the_altpll_0 <= internal_phasedone_from_the_altpll_0;
  --vhdl renameroo for output signals
  zs_addr_from_the_sdram_0 <= internal_zs_addr_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_ba_from_the_sdram_0 <= internal_zs_ba_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_cas_n_from_the_sdram_0 <= internal_zs_cas_n_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_cke_from_the_sdram_0 <= internal_zs_cke_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_cs_n_from_the_sdram_0 <= internal_zs_cs_n_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_dqm_from_the_sdram_0 <= internal_zs_dqm_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_ras_n_from_the_sdram_0 <= internal_zs_ras_n_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_we_n_from_the_sdram_0 <= internal_zs_we_n_from_the_sdram_0;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component nios2 is 
           port (
                 -- 1) global signals:
                    signal altpll_0_c0 : OUT STD_LOGIC;
                    signal altpll_0_c1_out : OUT STD_LOGIC;
                    signal clk_0 : IN STD_LOGIC;
                    signal processor_clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- the_altpll_0
                    signal locked_from_the_altpll_0 : OUT STD_LOGIC;
                    signal phasedone_from_the_altpll_0 : OUT STD_LOGIC;

                 -- the_cal_dac_code_pio
                    signal out_port_from_the_cal_dac_code_pio : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);

                 -- the_comparator_pio
                    signal in_port_to_the_comparator_pio : IN STD_LOGIC;

                 -- the_gen_code_strobe
                    signal out_port_from_the_gen_code_strobe : OUT STD_LOGIC;

                 -- the_gen_code_value_pio_0
                    signal out_port_from_the_gen_code_value_pio_0 : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);

                 -- the_gen_code_value_pio_1
                    signal out_port_from_the_gen_code_value_pio_1 : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);

                 -- the_latch_pio
                    signal out_port_from_the_latch_pio : OUT STD_LOGIC;

                 -- the_led_pio
                    signal out_port_from_the_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_mode_select
                    signal in_port_to_the_mode_select : IN STD_LOGIC_VECTOR (1 DOWNTO 0);

                 -- the_sample_and_hold_pio
                    signal out_port_from_the_sample_and_hold_pio : OUT STD_LOGIC;

                 -- the_sdram_0
                    signal zs_addr_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_cke_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_cs_n_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_dq_to_and_from_the_sdram_0 : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_we_n_from_the_sdram_0 : OUT STD_LOGIC;

                 -- the_switch_pio
                    signal out_port_from_the_switch_pio : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_usb_code_pio
                    signal out_port_from_the_usb_code_pio : OUT STD_LOGIC_VECTOR (20 DOWNTO 0)
                 );
end component nios2;

                signal altpll_0_c0 :  STD_LOGIC;
                signal altpll_0_c1_out :  STD_LOGIC;
                signal clk :  STD_LOGIC;
                signal clk_0 :  STD_LOGIC;
                signal in_port_to_the_comparator_pio :  STD_LOGIC;
                signal in_port_to_the_mode_select :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal locked_from_the_altpll_0 :  STD_LOGIC;
                signal nios2_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_0_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_clock_0_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_0_out_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_clock_10_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_10_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_11_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_11_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_12_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_12_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_13_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_13_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_14_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_14_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_15_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_15_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_16_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_16_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_17_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_17_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_18_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_18_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_1_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_1_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_1_out_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_clock_2_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_2_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_3_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_3_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_4_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_4_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_5_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_5_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_5_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_clock_6_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_6_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_7_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_7_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_8_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_8_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_clock_8_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_8_out_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal nios2_clock_9_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_clock_9_out_endofpacket :  STD_LOGIC;
                signal nios2_clock_9_out_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal out_port_from_the_cal_dac_code_pio :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal out_port_from_the_gen_code_strobe :  STD_LOGIC;
                signal out_port_from_the_gen_code_value_pio_0 :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal out_port_from_the_gen_code_value_pio_1 :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal out_port_from_the_latch_pio :  STD_LOGIC;
                signal out_port_from_the_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_sample_and_hold_pio :  STD_LOGIC;
                signal out_port_from_the_switch_pio :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal out_port_from_the_usb_code_pio :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal phasedone_from_the_altpll_0 :  STD_LOGIC;
                signal processor_clk :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal zs_addr_from_the_sdram_0 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal zs_ba_from_the_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_cas_n_from_the_sdram_0 :  STD_LOGIC;
                signal zs_cke_from_the_sdram_0 :  STD_LOGIC;
                signal zs_cs_n_from_the_sdram_0 :  STD_LOGIC;
                signal zs_dq_to_and_from_the_sdram_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal zs_dqm_from_the_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_ras_n_from_the_sdram_0 :  STD_LOGIC;
                signal zs_we_n_from_the_sdram_0 :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : nios2
    port map(
      altpll_0_c0 => altpll_0_c0,
      altpll_0_c1_out => altpll_0_c1_out,
      locked_from_the_altpll_0 => locked_from_the_altpll_0,
      out_port_from_the_cal_dac_code_pio => out_port_from_the_cal_dac_code_pio,
      out_port_from_the_gen_code_strobe => out_port_from_the_gen_code_strobe,
      out_port_from_the_gen_code_value_pio_0 => out_port_from_the_gen_code_value_pio_0,
      out_port_from_the_gen_code_value_pio_1 => out_port_from_the_gen_code_value_pio_1,
      out_port_from_the_latch_pio => out_port_from_the_latch_pio,
      out_port_from_the_led_pio => out_port_from_the_led_pio,
      out_port_from_the_sample_and_hold_pio => out_port_from_the_sample_and_hold_pio,
      out_port_from_the_switch_pio => out_port_from_the_switch_pio,
      out_port_from_the_usb_code_pio => out_port_from_the_usb_code_pio,
      phasedone_from_the_altpll_0 => phasedone_from_the_altpll_0,
      zs_addr_from_the_sdram_0 => zs_addr_from_the_sdram_0,
      zs_ba_from_the_sdram_0 => zs_ba_from_the_sdram_0,
      zs_cas_n_from_the_sdram_0 => zs_cas_n_from_the_sdram_0,
      zs_cke_from_the_sdram_0 => zs_cke_from_the_sdram_0,
      zs_cs_n_from_the_sdram_0 => zs_cs_n_from_the_sdram_0,
      zs_dq_to_and_from_the_sdram_0 => zs_dq_to_and_from_the_sdram_0,
      zs_dqm_from_the_sdram_0 => zs_dqm_from_the_sdram_0,
      zs_ras_n_from_the_sdram_0 => zs_ras_n_from_the_sdram_0,
      zs_we_n_from_the_sdram_0 => zs_we_n_from_the_sdram_0,
      clk_0 => clk_0,
      in_port_to_the_comparator_pio => in_port_to_the_comparator_pio,
      in_port_to_the_mode_select => in_port_to_the_mode_select,
      processor_clk => processor_clk,
      reset_n => reset_n
    );


  process
  begin
    clk_0 <= '0';
    loop
       wait for 10 ns;
       clk_0 <= not clk_0;
    end loop;
  end process;
  process
  begin
    processor_clk <= '0';
    loop
       wait for 5 ns;
       processor_clk <= not processor_clk;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
