��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�=�}A1��=1�<��xr7�n�?��;�MHc ��c��Ɨc�ɍ|�w1�ag�j�J�gDBʚ��n�N���a�� Zs��Gb��'�[����_��.#�2��*���|�PNž�0t��'�֩�X~!���i0��A��-�xI'O:1�T���v��W�r�� u���ڍ3�����G����Lֿ�^PQě��zg�nJ����*��EV�I�����u�杇�e,[��l��9Љ�`u6���4�
R�ox�uT\)F�^a�¦/��`ɁK�<��]Ñ�tt�GGe��[�]GO���Ŵ_Kb��f�Ok�i�(���\�,��br;ғD����1�Q������$7�N�����S?L��:�sJ}��%oy��������3�ڴ`��?�le�9��<m�P�y�!�!��sN�E��k�+h�602y�n�AtW�����V��N�"{�042'3����L��l�d���E�3�����Li�&3�����o�����Kk��:h�A�,:qoB�qU�g/�_a1hl���vo�$v����3��4�?-N[����w ���nG2ڻfod�<m�)�������h�x���n.��q��R��^�w5��76�� �8�m<�.U�@�:���i���jH��Ex�Ю���N����.�5p�V�l^�������Ft=֧@{�k;Ee�y�դ��K��Y%��b�ĸA;�QC:��������F��c�A��д�~I��O�,kL�S���q�eH�R����܅�g�2ۺW�M���?�!���;��b��\v|�d����^^�Ȱ�[��r;�e�WN��b���t�w���KĬ��O�y���-�gYդ����m�3�Fbպ����u�@�TE����Ȳ��#���I�>Dں�GgQ�`(��	� `������H�p���X��X��i9p�s��jCLa�'rg�_���ZǪ@��fͨ-�����Ia�a�i[�73����$��.�5��Y�׼2��KÒ�y����$��\�M�/�s��s��4�37��Q�%z�O;h�T_cD~�?���&���YfC��U�PJ.�?	�A�#���dm/�3G��Z7�o/!'ϐ1㘝g��,�P�t��K���w7րX�ȼ�~�����*���bQucv�����H��������:4�O8f9�<̠f]E}�.�̏4���B���;��H��ɫ�p��˭]�����'�eKR����E�"DQ8*�«���¼���+�ߖjv������V��hI/Q��ի��O�=�w��*}���q��Cq��IKL3��p����K!���d���iX#PP�Ź��4������������9�;vI-�C4�`���"�i��رW���H[���t0U-���gk.�<�����ZݦO���l�B�hd�#f����Q�ߑau|�Qg�6�P����.W�:F��%����X�)`.��:��e���Rt�;����õ�eНd���+�o͗r\�?Ծ����5\D�^��>�96J��Ȱ�3�bVW�NV\�}�-G	�qq2��m��.�?&���R�_|����W���*�`"����>� eF����"��o� q���	�i���s�B�@� IӴ����)��w��C��+rɥ�I�Ц�f<�����X�g]��S>�|bV��<{�VTGys�̣D�/�u�e�1S^k5�-
72�B�~���-o�Ed�u�{g��$r�n������I������Q�u��6���+� $�9O��j���h�v��>��{Kv�E¢ފ��H��^K�I�_��-k��1��?B��U8Y������	����z��ۅ�\oD�q��*L/�#a�Jh��m��3�sLg��߉D�e߀��s
̂	�H��H�,���n�t{������Lu7*����4Zx��xt0���=k�X����]�ML%��PqWV3&���G} 7gg���{櫫�*Y�lc��~��������:�U�ÁٽT����`�D9(�2N,�8�����lb�s�S8~��������-�Z6J}�tl'�P��qp��]��:�7�'��`��1U�i*�ӟ�	GCR���+���@����>��� &��!4�y4�w�?��	��S�-+䃠%�q����4��?tJȦUA�ߋ(�$�-2���Fr]nmR�`6S N�y3�¹��o���[�wm���>G�n���Q�x=� У�'�(���(��A�ڛM1DǮ��`]�y���oׂ�zSK�������=�`bٚ[؜i+D��7=������e��7�:Py� �d�#����l(�*�_�q{�|�qw��b��.�������2D8�^��L޲�d��d�gkK��i:��`.]gdV8t�v0O�UvU��$	[%��{?����^�>yj�?O���j5t��us���-���Q�l�y6jF2����8����=ϕ:yW������n]2��a�Û�g2D:�`��r������R��.O�K�]�4.�jX��#8m�wG��_h�z1CX5/ԉ"�R����ڼ��`V�ա�������#��`f>���\�@��Z�o�ۢ�ֿ�s�k��?=f�m�ZǇ��S�y����(2��m0�׬�<��ǂvV�M,�gk�xU��HF�-}ɓ2��f�B�W�����WLO/�D5{�60*��6a��K���PK��v�wB��^�첼?K�D;��:T�8"⣚���w�r�r��gJ�P���bw�Hq"���j�fr{�mf� X�wV+r��ܨ�Xg���l����*f�N#DOo���m!�KK>��C/����+R�ρ�Wl����)��SR9������`J+�N ��8�^a�Ch>�,'�Ƥ8h��!�2��J.�_½��,�ψ7)Ʀ�x��l�w�Ш�?n|È9�cp�O�D��m���7��V�i5������.�����+�}T��C5-�
*�m�V��`�;�)Zk�-? 	.�`[��	�踖�]p�Ub�7�C{�AC5<���� ~�|�� �/ؐ�|q׬�(����>��$"兌I�w�O�퉙��{7�Tw����~��X���os殜c�q�Yp��5�AA!<&�T$�2��Cg5�Ȭ��И�)���J8�:�E�q��u;�x~�*x�-���Z,1�W48�����&���H_W?�Ry�',���K&I����!Z���C�r��g��`A�:���w8���[�%>���]����.�(Щ����f6�$���,I���8,�հ/�I������U��9$^�NCc~�"�⦓���Cd�/�5�4D�"��oz����b�e.�ST7�7��V%��/������i[J��<��,W�9�@�J�y�"��gh���)1��E�U@B2���L���?�O\��m�S[�9Z*K��kl��=��^�U2FIJ|5!+��D0�X8��}�Y������T�K6�E ���ֲ�����A�~S\ү[َ�n��`���!�*F�&�e	������V�^CD|`���Pd��Nt��}���`m�77����Jd�V�U��TZh�����×�<�6�[�ߓ�"�c�G
�5T^Ye�1�2)Dh5�F\��� ����;��^'��ցъb+�O[�K��2��CQJ�c�A8��S ��N�y�+�H7p�H3��n!$��1!�&���e����E���|��$.�JϞG�l�iG�,<]/X���#�>UU���6|�T���V��5��z:�Cx������� SV��@(SC^��R�1y!K�Y� ��|6��I���h�:W
�Sͽ^Hw��%-"l�!..C4�fz�%��OB���>�<��r���a[k�\��G�����q8��Ur�6�yА�X�&�8�.�x��F�$�-Z�Eʏ/�q���?8�$�(BW측�s����$F?���W�&��rG���g��ΰ}I�+/�&�y+��izPra����H���f6&T!Xi��;C��x���Y<��6\$�K���s�]��-CXϐ���^r�Ph��Yb��T�+�� i�i�8vo���ri����cn�G�kI�µ�����_}�t-���`��S���Jq�|0���u�	Ow����E��;������~��l� �6�}UQ�
��՘�Faź��B4��7=�� ��j�� �8����F��e���ԗ�h��Di;�)���_w�S2��?ډ^����w*��qb���(K�NZ"�2��0�E��j0���������܏��g����	�8X�؋$���� >�?Lh�T�"!����_��Ghk�1�2����j�E�ԩ�C������D�'hǛ�T�u�C��k����^��B$��E˱���Mlt�e�Gqz\���}̜h�p�E�����^GZE"v���A����l��z���J��*'��MU�`E�-�8D}����ؘ�ہD��k��Md�s?V�rB��Xp�����l�&�,~�~O����;��" "g�ǒ�~����]U��}My�~���߾�%���ݽ���p+��?��(����{���ԬuIX��°[b��
֢�� R+�Of�����u͉��e�ȓ��^c�9�!�X����cY:*,��>�H��d��'�x�
��L/��	��v��P���f]�E�v��wa�=T�䲬��J5ڰ/�y���^R,´H�ʠ�HS~��BB&I�Q�*v!.����x38W]>�K�@������ܐ���G��r0P�x����8>	H����$"��fE6�I�: c)`Ij����j'=~��<әn�ꥤ�&v��kv���N�+��)ޜ3��c� �jk9d���=%�tc�7Xʥ3�`�����וIU���@/i$�w���uCd�� �tie�RF�&��֍�4�N�p��*��b�!�w���3q�G�	
!=��5!�x�Ŏ���?����(X���~�T�yDH۷�<�I��|��Ny�
�A�`)c4��ln�M�f[�y���P�г I����:�0�W�C� �-S��Sd�9��kb���4~m���MY��!���E��c�w���Wa��)��р��F"*�C�����jW��?;�ǒ[`��W�h�%�A�DwdA��? X5����?}�����&�����L۸Ida �Th>�#drd�9<<�x'B�W���)f��WwT�Z�#�.�!�q�&7�Ҟ�O������6M�̖D=�Bt�΍Y=�dXR�t�О�Zv�(V�
��x��V�gOHmb��uP�p.����6�Ϭ��Q�t�0���5O�
�_��"a���w�ױb��"�L%�G磝�;�22��k;��k���o��\@3�:H�8'bƩH��R��QQ�zX�оR7o�:�Zg)8�A�[+Q��#��u�11�,�c�q���ߐ��9f��c$�9:sߒ+q:ᕨ*e�-�8�8A��c��R�7�`��1"|��!uå7�����:�WV˿?ėN��Z����?>
��8*��Pϐ	q�8ֈ�N|įU)�0�oc{�u)[z�"�ְ5�nC���;K�n��ݬ���ɩ�PK�p�4)c`�6O�&�~�<�}��\�c����W�ΨV��m���'�<ZSl�;]�(N�� ���H��������,�)�̸��8	����bQHׁ�1v��x��6H$]6�1���M�[�b1�D(A�H���*����a{C����<M�#���+�4���`�e��g�[�����yA#jK@V���4��H�e�A�
���ۙX��l���ځ�a���k4N$����oq3�lk�\����Θ�IֵA�60���i�&�5��7�s�%Mt�df����d{��\^;y�[
�ګ-���J���A�Ϣa�vnNTRHZ�:����ز.��o��o	L1Z�6�[B���4�~&�lfa:�ʾ&��uSL'�Z���	�����yiZ�`�WZ�!A��=�g�|��<�����H�����(ʙ�� z�6AITe�qb�x�x��L�:�Xs4�͑O��C�MQ����p�����%�j9�g}/���P)��V���W߱W���c�ˋ�A�@ld[��|��@��Ժ;x��H*P�j �j��)�Ʀ�(�q���$DDy��P�-����j�x��օl�kM��:�v۽�F���̉��/]��9v���]T,��g���b��I�=��yoM(S��ZR�y�K�'܏lNT�#�.G���������'�@m�	���U�^��QE��PdVb1��z��8G���'�]�1��?bO�$q#ϒ(�PU�>Ř�w�I�HZ�f���_��ޜ�3��cu�k�W����ڡ",��DbH5Ә]����0'��g�Jl���L?���WˈP̦��z,Jb���펫�����gw2Y�q�����㨏���?�-sM��f�@k��/��n�5�������	ˁˊϵU�h��'��U�3�qzDeB��C� �wX��hu�^LG��ߦ��C^�(�m� �w��6���U��[ �ya�<y�>l�G�=0�gl��ڏ�IDs�K]
�T�"ŤȨ��x���ʆ5�,��'��� �$-�nK-��&e����v������\�����O)1�ʀ�g\�2�O`$(ϦZ�P00�r�y�ݡLkL{��K����n�w&�=+�{��b��6 K#�����D��U��Ʋ�r9�g�ˋ$�ʦ �ێ�2C��\S���\���; =H��EH�I�zA&�����!]�-����k�6f̜��r��ށ�^@�|=��Y���%-[	�.n(�F50K�6*��}q˓_�ȴ�a�hO%�� ��J�--��%7�7LX���r�[ov�����.q�/��}&�~8�di�,�J��B�J�
p��z���N��3
�Ѫ�AQ�;2��D"s�ʇ@�.��c�q�|Q�o��DJ$̍�l���Td���5�C)7E��	��oЇrMSG�r%�)A��9Z�݂��o�����Y�8�IpK�"��RЀ�ajf�Ή�r2R�/ך��� ~1J�E�%�9��e������7�d����+"_�G�"w�1j����L�
,R)_��Z�-��W~�c��(�QM~�A=7�c���%��m�.�:اn
!L��TE��p�i�o׵���\����Y 6O��TA����6о X._2�{;K"�P�,���o�u���s#	�n��Z���(���]�YE�a,�!��!3��$y_���-THzHf�I]�g�7�yw̳0�'W��xCw�#L��H��Hg�m�lJ߭�%��ɡ���w���f+�(z�;§��ZܸJ�e�ѫ�c[�?)�n��f������ݶ3�7���V����Mc�u��4T�����+�4fn��g�G#����#��]�x�p�2VwV�.�ݜi�;A�����^)�"�)O&�) ���mq-�}7{0���߇ ܩy����(Ӭ��5u�Q*���n�grH�-v��՞��(j��f�/w"�Ϋ� �
�4���5Ŀ���#Nk���d�y]�n'X�KHu@,[���*�4y�.9������6��iF�,�mn��$�iC��u��:&�g0��虑��!��Ox��>�.B�û󔭭��_��Z.��#z[LҹDL�ػ�6Y;�V>���_[}=}�g�Xb�������~!�h\%�1 V�<e�9O[���X/�Ru���KI�W9���MBT����!@���ۆ���x���O�����Ͻ�LP����S������\��p�� �hKHG�@�M枕��(˕߀����W�������.�0��sqy���ΠT�sZ�({����c3�6���~B��FGM�mG��b�x���55��n��Uf_���SF2�d-��`������G�QV��bB�����	�+��64����p�K9�⥝N-X�#KH����-Sw6gnQ>���S�����A�N|N��V�Wt���d�W��Ԇ9w� Fv��!>��%U�M��_n��@��]|��"� �h��;3T�K�� �΄{���Ue8�J�c�o��'�N�'-k:�Є�@��g�Y{�F��9/��gئu�t���.!?q8֦Ow��|���U�]�э-2�]\� S����3��>Ƙ눓:�_FiH��up�K��ؘ� �jped�� ��K�嵚v�A�ѵ��yH����v?ef,J�S(�km@���g��Z2��� �H�k�5ޒ9�7�~hf�q�>���=߷˄����/��=@>������뇧X�V���VћH��2��=��Mqҫ̓t������c5{��}��Jd��h�Ù B��ە7���*���{��4��2b�
�n��MfǄ�пr�e���S�m�Q�e�t��v۞��Bp�Jq�)��^iɺs�▬ډzvS�ǔTT��c�u���Ie��!_NDx c�����ݽ �>�ED��<�w���f�0��nH�H��0?4@	�;�d�a��B�$2���{�ns���0���u@���J.�I�W��d�f���!�ay��߄�m� M��;�I�M4(�lu���|�����H���K�3�Țb�y
�汇�z*������d��?n�5n�@wx�W!�;��H�S� Յk���`��w���zг�s��?k�<���ՎT�d"�6��"ߘ���Y�%� ����fL�}n�{�p=�� �flt�%!e܆M�O���d!�O���l��4帧����-s��m����,;�M[.d�f~V1��nI��+����|=e��&c�׉��=tT�թض�x��T�{.%���
@���-V�Ӫxc� ��(Չ��F��y���&rEс� ���Z��sSg��ѣ��lI�+���킄�����Hu��#�y�ѵ@�-������M#�☡�&��=�oh�R���$O�����Ɨp��1&S��G���+��A���G�SR
�%Y~K̺%l�w�؂��G܊��\U��E�]���G��M�-R�%#�>b7L�C��P�U��㸢Zuo��4q�^��U��mL��JI?W:�1��
�z�Į��`����6��J}ק}�^��w�T��U?Wl�J͈ȹ�=1�z.S�#o�f���˙��I�x�S"��@�d#/$���?p��pf�1����캩����x��^i�mA��,��t_*��x)��u�ʲiG��470�p>S��54�FxH+�WPJ����0�eTӑ�����a�D�ᗭ��_�j�:�ULPue�Xl�������vc&rm�m0�ay;X�]i-����4&�ao1h�H*��1��?'Ѵї��n�P�B�!t�Z�ē��pk��Bʫ]���:���� �l�F�F�*N��C.ܐ>I�'�#ѱ���hL ��pW��;��e��z�/G�T���RN7��V}o�۰�3���sf1�A�8��!��GLH�u?9 P�U�e�%�"l�f�V_�A!|����c�����đ�=%xq���A~�I�{�����7"�+�w�g�9%C#I�U��G�8[���)��f�ߔs9�)ad��3f��<�fe����[�f���nGQ_�Bp;�)��ǂ���=ф�$c8�xp�y�����"~���5�*%���I��7"����_L���G����=�D��	��0%�K����O�02_���O�Q��$�/�e��_S��֮,��%�P:��5�}���x׵�@B�?�c�s�_{fub�8S	�!k7_��h&�ђ��<��_i~�莾��?|/�
l�����7u����!m�q�yޫMs]�y!PB	�]����)����7귡�J���6q�7��L�A�Jg��Ǘ�ֲ-�4��q��S��{HY,U�B`n٤J�d��呤Y����Sb��T����7�#N��[�HW?�U��竄�J��bw^F��a�X�!i �i�"ߐ	����B������똈b��J���t�C?��!�@�[��q�X��m��.��.⟧�z��U�����%�I^��T�H)�+�W~K�%��d�NGK�Ā (�c�N1��)���d*g� (�j�Ì�́�Ѻr/� ��&柍EW�3�:G�ycL^�u�m���A5�4o���X�e6aZ�DH
x%;�C���1ƚ� ��k�@��<4�R�������+��s��/��
 �ƩIs���V¡�]����oA���ߊ����_l�-���	�B�?tb�.��-���Z�A�!���U�"� �+�U��șLf���jDFGh�_��6���s�*C���L�u!n�֤߷c4&��o��н�����fe��g�)-4%!��	�������a�%���i� �rO��}��den��g�'�
 ��Uu��rR�X�~��r?��5�<�8�^�w�j'�����3��JxG��1i�I����!Q2��Φa=:��m��̏څ�<BT4	���������$��0m�o�#��7&n�9!���@�-ޜ��H�ro9v����l�aF*^.�Z�{�q�v?�e5	4��IqTi�`@���
6P@�������ف���[o����
��S���[]�7%L+h�u��3�g�b`ҏ u���QT΍G�ו�_y����7����m�q��N �4
�R���5�����I�$��-��nnS�'@=�Q���"����Ym�zuǾ����c��=����];93����?�����B��R@:<~�.�;���"-z�y4����zDu�Z�ǩ��/���>����r��-i!�)��H�� �ԍZ�Ddm�7s�<�Í)D��Aͫz\�����4*��^�[WA �>��	���k �T�IalŌW��:���&S~��1����I<On���<�g���C1{٬�)n��3N(�/c�o��
 ��=��s���<��	�+�~	"l�~�=�� ����&@g��;@�ħ�sg�R3����OR$�I����Ͷ>|9l��L��1啕�+H���x4�J*ml �y�mP�@���=1e4d�9�^ُ\���V#�yr}W��C\�I!�j?���b��)EH���҆nN"4��t��dr�P�N�%Dl�=�+��S�k�+N�d��+�5ina�2�S{K�*q�Ƽ����l�����N�4�^'r������-��$_�
�/�n����g��\U/T�����s0��Y�VɿkX/:��aDmy�ˁ��^�jt=9p(��\@q��w�E�V�/Bj�	e��(U@ᝲ�qM�ddΰ�ū0黎mi����
�Enr
(\�Ӯs\�u'H���Σ�XC��aJaKuD�Ǐ6C4�W��u�c`�3�ֶ3�.���O{H�XW�:�[n*���bw��o:91���Ce�]ǂ�XV�w(�@�^r�a�-�����7���F� _:�hC�G���	.����I�&����i��*�j�1����ڑ̤�5��'���m��]6O�NxƄߔA�^5:ױ�\%��1�E)�<�ͦr�>7d�E<��-r:� #�qէ$A�26�,dM+����u_^�S��Qzi�\x&�������;��]�̞X\KF��=o���c�־팏���?�{j2uKz���[+�I�N���D�bQQR��٥yFMy��ކ���g�������z�j�Q+m��Zk�Ӷ�s��E%{Pv�I@��8Z�!۬!�~oa�!b ����0K���/C�d.��fǞ���܁�Vy�+c/�š�H�<�8k��9��Ȼ�	~����T��}�D�Y���ZH�ؐ*U��)�x���B�À#Ɲ�%�'����,�{��gC�re��Sj�Z��B���,ST{�	��-��A���zx��'�:7��x�� ���/����� &~b����] h?;������6Yo�
E( �Ѫ��ñBp���Ц,�i�Q��d���:�@���W1MϢ��
��� ���涔##P�\;f���k�F��}������F`�ڧ)��C"���p�5�ρ+b��*8���6Xw%I�v��p?*��dFY������Rr�:Bc�i
�8^_7(����U�ܶ���h}����-] �X���e�i�����]�)n�8S�b�q�����GG.WƤZ�)��)~��	?|���K�s�+�9Z�Tڻ-�gt"*���z$Ԣ-X)�|!AA��:c��;�B�O�@|6C��
<�o��u�m�������J��o��Fa��� o�S��J�a�a0-bZ�$�預/Y����hZέ�^�qJFe��j��a6�n*N��}�z3=ȝ:U��W�u��F�o���)[�CCr��t*���s�4㣱�ւEw��+&��`&�g��Z���6�����~Y.�{�H�	7��,�Y
�q�~-,�@������Z��gY�ǚHd�[҈ܸ߭�{M���OXP 2�*�ӳ�*4$(�(p�P�:��O��I�Y�[��҅� ��|��
����乨Zd?P��4��Ư�ʷ�����|��#��`�xa��Nle5ix�'�7�p�=�lb��lث-b�g��7&���@#����`�,�蹖ɀ6��.�w0A����Kv��jU|ZVT`�����8�����dz�c���(6���i��5Q��Uѻ�k2���.����4��B�}��Dzil���a�d�������Ùh�b��r3�(z�l"�h���}�/��w)�f�����&�B�j�#$�56���2S�~|�R��_�;�.C�w��tY sJV]2�O�K3k6ɢ��2d�����l8����v�H@ys�X��\��7��j�a��7��ɞZ��`q�����p0i�?4_�?��=���&�Q�`��x����^����u��]aXHw���DU�����r�˳�yU��f��X4x#Fp\5�*��҈L;��SߚH�,O~��^��Sx,�|�3���ߒ�#"\�K|+��ݮ��\!���"�	F`Xߥk�l�1*��dZ�땲�LMN�L��/�F��v����@?�`�7�+�"
R�}����3�-��S�c�0'�Tx��1;�!1
���(���^ψK��cC� ���U�gq�D'� �hbA7��/�D;�� *������q�r�	-ͷg<�VLf� }�uM�-���-�Exr����0�ύ��}P����Y��'/���a�l*^��O��0
�'�8$�����|`��v�l����V3�+U�T�~�^;�7-�G�s��uU�b�L|R�5qt�����Ot�{.jp�݇'���C��.4�j|���]�0|ik�����P`�ePx�݌�B�G�d6��� T']���kp�/���E�9�&}���F�h��Ts�.U��[�?��f���i�G�Jx��
.��O�_P5@�q/�>u��&/q��D�^�0�&cN��z�6�W�=���d�-��"b�eY�����M���U��m�P>}�d}zt-^r�Ś�w\�A#�Pck=�ч3eR���D��a^���[*�01]�f���S�K�o.��櫡���
��1�:��V����i9�a)�����ۘ�����&N����Sf��?ކR�ɉQo�%{�l�g�9G%���
9�Ժ�7�l�C�_�>c�S���T�"����L���#��0�vے$&%��)�����`�i��)1Ǥ��c���B�B�r ��;;nY�A��B�<DJ��Qb
�,>g���9y�+�א��Z}��t=a�ܽPA}g��hQ�3.xa,`�s���R5үWv�_�S�Q����G�3q]���|R}�ހ
�wRS3��{��>7�Mt��	HD��`�Ds�#����<��&�͏69�2v��3�z�YF,yHn�*�d�z[��8|g%��e��	��(�/�����8�JM)���pZL^0D���jMPi>:�aw>�0�,
�_���G�]l[���Da��v��
BM����ug+M7ɂ+�[������D'Nf?bEb��HU��<�
�s��{�	c�;�����M��p/j�d-�:F�HNx^��U6�T�s���gӉ��r����/��R�`@�������/�۔g7�B1�L�S���L�-��@�����"���-����{�4z��E��S-��©Z��kC�F;ؿ4f���i?X?�hH�c,�EpMw�c�\I�*͡�Q�6�����q�th�N���ɇ�P�x�h��D�H���P ���	62��@)�ъ�a��}og�>��l�dV�^�����X�ߩ.�c'%7�nƃ��C�|$��::���&��v�5�5������
�Q�2&�˥�bo����XT. �� "�O��WjO��D.7��1� s�|K�@�����z���J+�nr�Y�@��r�@bV�7�%8�O�S&��WF��b�֚T��: �R���fc�����p:�dL�q�jXG��1������27g�Z���3�r~�I�WZ֝jma���e~A�X���_J�^K���3���g������a.4�=�z~q�c}�s�@��ŝ"�{C�Qq�+@U���:��+���zQJ�l]��;�\���ܳ�3 ~��3���'dX�uM��*}��k���n*�L��4F��r) 8���?\����Ǽ�[��	Ч�m~��4���DL�V]Mzm]�!��~|Y���5�xI�%��n��%��L֖S�mV�v�|��29�"7��kU�Kꓳ��n�!��~
`���y�ؐ)Gخ�,�!���p�}��У���!�3�<z�	�T���t�F��|��H�V{���(h]�t��[܋Xj�4�Ryų �bB ��E ���m�
�l�|����#��A�/�E�����m�A�  �^�2s@eR��̗�x�k�M��Q?$�8F�6p�LZ��y,k9N�Β��K��,�'��fPg�$;�⪘4�
һ�� ���j�k����iz����
����v�=��AE�P����f��3��q��.�0?%�~¢��]k��<�*����t�cj�2��a�T�M�Ӄ�3n��QR��-{�G�QhLK�6r������Q��U�n��ҲK�D@/��௤�/';d��N|um����) .{lU�9�b�~�>�C�SFCO/}��K7ґ!W��.����b�7=�rv����J:�ˬ�U�����D����.�<��Nn�=ǛLb�[V�s�X�y������
�V9D���#�>���7�<n��^�M�&����2_]p���<hltvhw�l�(�eT�7@G���K~�ezK[nKn
��g����.Qc��� �- f��>�7&CC�����Gpo� ���Ȱ�qib��׀-8�eC�o�Os��G���Z��x�ҥs��!��:t�Ւ����.������M_� ���xZ3���]���dn�=�wBw����~E�~ ���Ѥ(z�.�ãF�M��g|�+A���JZF^6��@O���1%���1!&6;����d�h Qܘm6F�T�R[.u��~w�1�\ݾosO;�%�HVhd��*�����n��'�CK���O��4��|"G�_�A7/Ѱ��n��@�ōj�=ϔm�1 �T7�KY�Ī_Y��K3T�_H���&��K������L�E��6+���r��F�ytHlE�ģ�PLi׊|��N:9i��g��1"����4u4w���S.Jdz� Q�����Z���]�;�E�w�P��|��0�I2���(�ϕL�x�=�u�'V���a+��z��aԠ��"��Vķ��ʚS�W��a㌀��	=�!�#�Dg�N�ɅoN�"��PrC��+�.�:��s�D[J�i��4l�Kq��lv�!���7� �-�8],[XF�NO`��[$tt��%�~2�^�5e�k*-l1�I���=ϱd�µwT�y���f�v��r�ق��)�O��b7�if��7����ɣI�4��qrS�"=�V��7!�ƤZ���aÆ�CR��0�$qKʯK���NV�3������aF'S���$��B��:j���1���8{Kt<���e�21������p�Wa^��;nAiX��WN�6�jږP#��^���
a?�y7R`u]��'p�+�嵳e�k0������c�.��9M��G�~4�� 8��p'�oP>�����n�؞O��%u����܆�]����{"��D�?���%�*@v�Ͳ|��E��v�U�w�D���f�4�x譻�lJ�WγߚVҞ4���wB5����Q/+�I.�L��#*� +B=!t�49%�J��T�THF!��c�v��|&A�͙�b8}�Oo�?YAN�X���»�K��~��ky���f�"p&>2�� �����b�IDW�z�y~���g�]�Px��	(�~,/�j�8��ACV��%�W����s�T��!�:��L!�:���}4��4!�����2��6��q&~�,�B�[��	�Xh)���H�>���_5��\H��BX�l��?��"k�T��)������-,[,@�t���.Pۀ��W
A=�,J�ԍ���YF�9�-uAc�O��֟Ӭ#&���РT|�"�ure���ӷ�x���O��+��b_�H�O^/��r��}Yd��=$IɷA�Sx��2%[#�q
a���;����ǧY�wK��©�I�#E¥F!��{66�/#�Wv�h1|���(pG՚	��-�W���x�^d|��;��ެ<�>�W�M@���Ж���cEe"�����*c�r��Dk��=������]�"3���N�G�'����^��+��lO��z:!�*$��O7���Y$��v��nt ���&?�b*Ж���6n�ἔ��(�����ưCc׸�5��O?c!�4��b*M�5o�<�O�=7���;�*��2jO��bс��V��x?'�)�yIY*e�_$�q2Gw�-|+	�����ů"�3��#�%�'LW⅄�[4� �:��®�aO�a���ʴ�}��Hu@��DǋRt<�>Mw{�{�b�
�|����ҋ�T��7���S����VE�V�7$�U\cm<1�G��u��Xu���\A�� F�)]��o�>�1�lU�t��|%.��k��j�Zp����lߠI?z��<ò�웝��;Q�
�;�C��F�����F�B�*Q ����PA�H�I<26@ދ��fJ��V>��6�V���J��p��23�����|#	�<��Q��Jey�B!EL'Z)��?Loj��m6ȍ�=�����)E�(�c�p�Ԯ�U������Q�)'ɪzxy��C��M��Kܽt�^DU0��ۂ�}��Z�C�y��%6�k�5�A6�͘8Ȯ4]�Uvk#�j��pc��$�t���R"�gpvӂ��[�J²qH��-@��M"��0�c];�Ko �3~��D+�^kJ��=�;��zGor��&�b��qη�$�>����7��fp������^+��Q��Cu��=H&q�t~M>����#'��Z��̵݂rl�DB�BE.�L�!�e�4dE�1X.�W��V�Wd��kdu X�)��?x(��Ш���gtњ�HJ��E���;�L�e���E.]�:v�G�M9V藄��+)]�������#D�,L���mҍ.�j��L�3�����VV���	�J ��6���LCO��X��8�`���x�u���&���/ΐ�%u�H�� ��p�Oq�+�����p�g�{���[Q�Ws���/�yBq@�H��k�Kp�~����d�9~#��Ԯ��	�F�g���:J�UO㌸���qH���qfR���WwE��&�āee A���19��@��<�˚@��M�����o:� Ǖ]�k���i����̹Fܤ�3IV�oЮ�F�~f��<t�j�H
�iC9~���O�L��&)CH6��}�[�Q�џС~�8�"�t8��q#F(�BuE��xT`XS}��'<'P��\��:�����{]�q�S��l�t75��	�20���Ӥ�`�0�[�g�r���$�s	�$���W��'�ʈ��=f�̹�VF5�I�8��K����  �$6x�j�jer[�U���\g8a�G�0��I�c��}�C�g*;�َ���'�Y5��ֈ驵���u2#s;����#���9�g�).4�!X}�TZ�GV�͇wX�%��4~�.�߈�{�N���`?�E�~x��
�!@ǉV%��pE,S=�:(�x�\�2�$���i��p�S��Z�Ōj���Z�jsf��a�у�>�å��g_�>edHW��s��{�5��/��pB[��C���ވ���r�^���ů��{o,;�yn��|o�>e�/�E�şM򃇴��	�K4*�4���_�����J�[��'� d��p�E��ÙͲ�s�b���r6]����͌DY�
KfPmw 72�}�Hv��w��Ψ��L�S���-hU���𮶪���������X(�f���	�z��b������xw���L`��U�8���e���;}[O$��ݕGV�S�FE=)����/*(ٛ!���w�Me}񟹊N,@$����(_��nR�;�CTuOLxxH 	ܚ��dZ���D�����8: ��D�<,47!��%��6��������q%�Lw5�Qn>n�BTR#x�#W�z�V��&����H��(~�0���QmPo�48	K�l>7���\bٷ�T��u����$S*��B����VP����'F�EȎ��C���z�X�@��	i�9��O7�ÙKX������q,]Y�޻�jyqt�$��H��᝛�ϴ�H�N%��P�� ����7���q�VFM�	p��|���Ht@�C �	)�:��(�u}��)�8 ����Z���)k.�u�����U�A�zЧ@cBJ���п��@m��8�E���!WK��Ku��2D���ӽ�uy� �%i�}���%2D�#��ɹ�ت�	L����B1�-do@9"�j�{V!�<! 4%�����W��&ݻC�W��2���;�q��kӱ7�Qtfa�����l2�ނUC�<�+���Ow+:��EB���Ⱈ��/F�3�G�n�� ���L����Cʑ�v��j�K�J�μ6�e+�	*�}�ȭڟm�o��e��h��l�ad[b���$�t��I"���v-\X�8�6o�@�Z�V�#�b̭��	-���iAj��]kӯ���P�W@���$���c�Rp���>.-B�UB9����|���7��g�g�|�9�IGQ�LH�Ҝ6��Q̞ƨ7�|��݆Y�<z_���0�,�()�a�2MĬyL�fGcξ�r��z���f,V>SFD׳
�oIz��"wj�yj�l���'��3��ɝ=��څ�՞�$�<;�(ں9\���WAO\��f�{4�Db���� �p	.s�aS� �����bп|=̯�U�^��L�ϻ�.��cFJ��b��Z����Ɏ�7�����{uY¿�Y�U��3x�ӊ�d�u#�l��샫{�X��8�9J�e.Sr�Jˇ�e��0�A�% ��ʩ�o��*jAmZr�`�,��D�桲�K��|Ӳ���	���@Es8��r
�"��::��eDW~1ݜ��D��<�B���1b�4�?�UϨ3���Z<�+� N����咙$�u��?�dЍ��KU)��[��O}ȞɜrȒ�\-�s +�iM���&�D�;�_�r�JU,o��'(�{���n�/숽�h�nO�ͮ#��/��ڈ��L���e�6(�����\�e����e��'�x�_u��1G��sܵ����ͽc�&1��F�O�_W9i�cL��~t ��������iV���'�j�Tn
��������=�l�3-��O��H�^ΓcR����]�s�=w8� �"�=@3>s=@N�"�t�6⑝b_V�ڨ|h���s��7� ����țe�5�������OdKGK����S-*-e����?���j?������t�\k�-�E\�Oޞ9b��|�Ә�f��-�3a�'�^#>0�v�'���$�q� sFߤ�S����C=�rt���:o��5�C���
�]�"�B�P�TK���k�Bt	4��g��2�����խ@�'�q^�a��'Ę���`���I�=�����Gң�5�/���PR����$�i��P��쵏Ϧ�&+�"jQ�B��4���l�=���KzL�U�ts���>b��Жꏘ-��o���[3n&}湺��g�z�M M�9��?ѳ�L�����Hâ���-}RT�[P?6Ʌ^�,��E0�7�s�W�����sL줜 ����+�kL$�%ZR��O����P���(Vr(���F�~�'����&��.ó��,� �%��<�_p�%��U><f0�u^CS�s\qUG�-�3�:����$O�M*Te�i]�p�eQ��)��[�G�7��G�f��l,�jp����C_��6�=Ж�]�Z�W��;乼������őU��8����M,1�#yA넘i�S��&e 3^7�5	�������8ZZ��ή,�Y�(�b@��M_��YQQ[�ny�׾�i�_�wP._PB�Z�����L���m�;�Ux%[�|�t���8g~ }��>����n����v0�����M��tY-!�i6�%i�>����*�o�D'k+���A�U�;4Z���7̱��/���	&�ͪ�eps�	\��{�Bv�xXK�ԝ�s�U����kg��~�6i�@(C%z�"�Yf�=T
^�pSj��k���S�i:������x�3M+����~Pz�4�`g���J7 �_y+�R����*� �kt'p �?Sx��Xu���?/ʖ�����UX���O��Q�6�� 
Z@v=O��/�lK͖w�T�����nEw_�h3Cx/�='M~R����R�7j�"�H�#�amws\TP�#[�R���	�jS?�ɤ�y,y���E"�:�t�L�	%0��X�u��̀�g�ڏ5v���\�^��s����ɉH��/��O�We��h�psvo�dם��؛���.D�K/�����\� ���C-��]K�
l�l�ox�ޢI���r@�3��{���3�]P�Cҷq��wC��b�4զ�Q2�c�a*ᦇ�A�hmO��\��"�U�x�Vߏ��|ѫ�l_D�["_!0z%�l)��ە�����l�L�&�&�=�X F��e�vUr�=��LA�Hy 8���s�Z�r��R���y���.p��"��I;�V�\��8��	.�-�MȞo�_X,��|T���ξ��Y�Z�:h/-��n��V��Τ�-�VF�,�hV�쉝K��\�h�I���-� Uo����7ɸ�#(����t鈫��A�< V5�`�0�C����v=��X*h�Su��~@s]s�W�lo�<�l�T5Gt+��G�� �%�b+a"�DT)7D�Ħ����Gk�8WLlB#*�""O���o@�D�5UZb�M���
�-v-�51�i���q.c���b�mɣ�eI#�c�A��`(��Įc=>0N�<E�]'Q�O8���h��[��vtL�j2���-&5Ll�WW�1�׺O�+gE��ޱǧ.lp�Y��#m���$��f���%��^����L��J�!qPE�H�JJr���R��Ǭ
�vu۱��	d��U=@��wUwO�FC�pI�m�׀�f��R�ԏ�jiZN��en6�?�)����gL��>�n�ֻ���6=Gu^1V��ut,g/bL���SV�&'! !A�z+��r��A���̜�I����74�C�}��`S�6� C�*9\A=_~�(=c�~�.m��>����~�斁���o�R��^g%ȩZ߬r�[^K�q���h�6�8�@�E���`9��J�[�kg�_��-������S�^D�8���S�٫AZ�1���a�#��.i�gq�X�H�*Gx���j���j�aŻBK�O͚�?}IˮR�@7���A�P� �&����u���p��lwB�+���x�e��@RDC�7X�����@����˵�D!��y��iwsO5o��ĭ#�p�:�U�M���e��qC�ٍcR��q�����B�_��3�nX��y}-M�9���{�$�E��]�p�?����c~!bC��Z�w��'���[\ar�8 ���%|�l׾V���Qo2'H���'Zʧ{A�ؔW��_t���&Á\� �%��T��Z�c��N��^"�1e�ŏ̳,E(t_�Lb�!v�Ɯ�;�����'��U�{�e����-�8R8@��d��K�,��ӝ��L6g/2/QBT�t�ޞ���ab�'q��t��,�e�7�5m&�<Qf�d�v�pT�?>T�U���fZ�9��.���)�o	�1�+�,��1yݓb����
���u�k��x�lk{J��G,3����7ɲ� �����]!"8Dn��A)u��`f(mm<�M"<�c'�ޫpAV��Uy��ಞ2'i����]
W���o��"�$�>��z!&�1���5�&���O&5Q��t �4 h�)��枆�*l��v�8FL���!�<����.<4�N��TOKk�K�����{�|�I-�S���C�Nğ���R"��Vu�nؽj ��,x��!4N�" �x�,W��-���8ď��%u䃂���Ќ^��z��� �~���0!˾��H *��$7J�-��W��lb�&K�h��%�eS��Q�FO\΃�k����1��B�B�R/��0H����",�,&^�
Εno�yRdj-Bst�4BQM��;��T��{�Vo�I�@��9�l���w��W�����a��(����l��񚒇������A���z�aZ�S��g����oh��!� ԏR��7�{�=��#8a�r��V��8�_#z��!�@�Y�2�TD��Z��t���L �(��9�&fT=�ī����6�V ��X�b�H��]_��ł]FD}�5��J5�8yт�?;Ɔ�K�4h�~[�>�˿��DX����
��Я�c=+YN�W��{^�t-Z��Ӄ�&� �w�$/ND��o{�PEs-̰-\1Ԇ��\=�(���=õ�(t鎩Z�[��$Zg�tu�E��1E��Y-�Dz�g�����"����)�}Yzs��ک664��R�}<C-pݬJ	1-|	0&�el�-��πs�y����"(�����f���q�ԗ���y+@GP�jËa��� ;u��XU��b��qɽ��2�o���8��IԂ�h�_Q#��ْ�%H>��k?�r#tL�\�c�ض������+��h�Dﱨ1J �k3�28#�H䣂��Ԩ	�\4Q`�o�����ՠ����%.�6&�{>������e\�U�i��Zʯ��2�Ѣ�ԫF��9%kaх �� ���Xwh�2�؊:�q�<�,��۽���P*ē��ęж?�@6�e�PIr�O{�� OZ�L#	��b���ӵ�����S����G��n肦s�,r���_���:�Y��^z��I�
�Y���<|�Ӳ�=KPF,�+����E$�a��ڪ���Y���,������Ƕ��_-��)���z���^��PW��L)_n5��g��B���&Y�&AY��Re��"n��Iw�n�x$vN�3�D�Od��DR�%���U�5�{�A4�4��dF~�̠ս[e�؍O�B7|���n�@�� u�bbn>�}��=�ͮ ,��;�F�C^5:n���0�x�Nk}l����nʐZ��A�m�O$��ډ�F5/�����⻁[�|*�m�� ����ߧ,覺ٻ��ƻ���`S�&qp�O�����5�����K�T�3@���w��-�����+fBz��<ELܹ�i�Ң����Jg�)�x�<��!J��خsߐ=�`��,�;4�wB�0h�K1"2x�}�<��ݪ-wL	+z��-���i��u����8��Ӵ�@T�Zz1+J/��݇䪳{FOcc�p�*3��'�#�����4{���{b�~�����b��%Ɩ���Q�?�4]\��~�U��%���-���&��+�nVnƮa�"O�ɨ��8�C�!I+$�M�Pd�C�n�-�s��@:6>�ϑ�z����v���A�w��x���wWv���r�6J�U��2�pf8��W\U>��A�٣h�Ʉok��am���
" )�
�^9]+�myY�m]�ŧ��c�Y+����T�RA3;Tt
�c��Ȧ׀����;��QY��V�ъs����X"���7��e�U��5��(�p�V*;���ş����W����CYT��68(��1���.rQ�k9D��߰���B���gX��i�S|A�@�ʚ�q�J�Zҟ�]�$���pP���-�4g9��p��D��҅9�������"�W8uP�!�|)ՙ!`r�2�F�����2S��,^0�K����s>�#r�D��oV���m�u]� Y��5�WPf�p:6��
}caBw���}?���w]\�x��H�cO���n�=�9i8�q���'�W�L�C$�z� �$~/(́8�r�@��C�XB�5��Su�t���
�ޤ�̝M퍱����
a��8mD�߉!��5|?�Î�eQZ�;�M���������c5ϕ3UH�3�X+yYe���
��8S��PÝ�+4 <���GQ� 5��x<�r��'j�G���^�6�f�3����|'�D؟�$H+����ÆN0�Vn&�'Ǘ���%��%������Rw�!�����s���q������$>C��B�9>�"���ƈ1�ِِy�&/�n�98�!�L���j 7��94?�@Q�^Eyq�P�����Z؛��I6�ڛ�[ʢt&h:�!����Ir++��t�����<�It<BOWcXw�Y鄛�w4�����_E/T�m���͗�D3M�X�	�`"۾�8DŃ��g��kZ��Sԫ��C�i
�D�$3��F��4b��Z|��!����$�r�W�G
�a٥�V��5o±�D !12g�&�G� ���	π'��'���B��}ĥ��휅��ٍ��*MI&oVs4�����0�+���b�������8��6;w
2!t�`]���5^���u�O��#������`��LqW��x��S0�{��'�T��u�:1�����M�*ϟ��1��2�Z��c�;:C �@�b�Ď���I�^�\��~.�V�i'Ý�C��S̪֍�Y)��(��^GE���>��@�3�OԗuV'K�LR�+FGal��'�R����G��������i�L���c,���'���<�b�ۼQI�N	\7V���b(���]��=��U�%���<Eň8��~� b-c������`�o��ya�����*�/�]�����n������~硉`�v���)�[�]c?��kU�b=���*�+���BN�t�U��	'i��g�p�����LK)��X�ԠT�(	9�+�`��ˢ6Z7��̂��Y��uP�C��̍g����7b��N- *���a7@r���n�a8Ti.��(T�k��$}����^1�ſ���Ha�6!!��=Xj���e�Z*��^ �w��xW����U��t��}�L���+�/?^m�aU�]��">ۭF���ڃD�S�{�*K�����x��	4�v�4Ϫ�F
i/��箜2O��-�&�y6��F��B�dm}O�H����av4�~�h��eo�:��8,�8�n_�@
a�^��-���T�����^�6�w|VyK^aI���%81L��6b�y�D#�-�ؙN!�����JD|4���8Y��KO��m%�Y���w%;���b���C��C����&�~gTNJ��ozܸ��m.��~!xi�!�4�S��e))���ɔ敔8+9�x����L��;~S!��T�)�3��	3}����@�Ve1(��w����wA���3��=� *�VW䱃#��Q�o�Pְ�V�Oh�ܯf%�� ���T	3 ���e��A���*)�G�,��.$�$BtF�F������f`�5�����g�/$c2��IMʰ{ښY��*2a���v�F��a�����&;�,o�-��\-�T���g����3 %��.ZR�ǜe�c���E-��ߑ�L_� �0 �m�B������Qe�fU�OQ욣%��=�fŋ�W� II�Uh�3��N���pzjvyq'�N��Ŵ���l����E��&�W[�~_�
?��@�U$��Gp#n���xT�)�b�{̗�v��ܟ�+�nV��콩~zA'UDgF�b��@'JJ�z��K 5D�Loȣ�^���^�P�.��Ⱦ��2��E{}4�l�zO��i_���R�u��~�f7�Ӊy�4��.;y�G���.�;<Ѕ��g�~1I8J�(��T���fK(�Ё*���w���;���8;�3ټM����M��m���XO����̶��/C�z�#���
�)���H��4!@����SŨXI@Kˎa�Y�%������<��r�2��N�{���&F,�f�q1�ʫa~�$o�:q�3�O���W�4]�I:ޑ]�c�E���M�t�fb��r#D�a8������X�pjb ?�qg���u��k4Q���^���$CF��*4)�AX��L�@������
�:j�⪰j~@�+p.
��U��*\Z�̽{����묓i��C�7�]$���k(2�2�}�˄�C�3d�����l�J��v������P�T���?��ܝ,ˡ�n�je�_܁\�������(ȫk4"I�I�D�<�!�e��:���]2x��h��ط����.�P��n�6�1ʥ(�U(�3�-%����X�
�m��IDJ��DQhZ�:�Ԗ�Z<�̭���_�ѧ��6N��hvĤ
�Kmŋ��]|���i�IA�������/B�g�U7r{�g�o�K���8#f,��L �
:��PJ�Σ��of���'U�,D*jLh�K�;�+�T[f�a�xh�Q�`ݏl40�0���WI�.�b�A�m��0V-�z.� ��x�*ei��f>�<{��[��Ap��iؤ�}֊Cm*#����-��.<P&��o��4�$0����(J����|YE���5Pꈞ[2�*��w�{��}�j��cr�Gm�~������Y�QVM�I%�4�޷�d�fZ�0>0��p��s6����a�rm��zZ��4aw��_U2�a���o�|$ğ���I�$ ��;��H�;4)�Sd��"*�J�W$-d���_��0��I��p�_�P�����i��1�%G�n5$��{�CeI�:Q2�"-�7�c���*r�����AR������Bj<i)Ny�2��v�%�V��[��fm����D�9$�Pl�Md3�h% |�m��CM�6�s�g���[J��t��a��2ߊ*U�#y�]�fk���	?�J�!i��걡�8�;�#�N�3k���[�,9�$ᵥ�ROo��]�4���U^,��}Cr�����Zp���̰�E�>Y78c�Gc ��F)�U4���7,��c	F:�$�4���.���U�aX�	ޅ��[���Es��v���F��\��krY�o�#l�q/��qD1�7:�c���
�3e� ��vq��}W�Z&-΃,/����
DG��䔺�Pw�&��vH�ۛ`J�~�A<u�.w];їd�?9oa����;��*mnZ�z��<v�."GV�C�5^|4vm�ˤ���nݮ�X�Z*Ng
���6�cB�k�^c��TjP��go���,t���zupiK��a]*�78O�'cXo�v���YkUª�(��x��R���Ms7�ǣC\�7f�e�GoXCU��ǼRn;�5Ϣ]�A���U#����X|*A4�����ט��ףN�������,����8h:,�H�%����6=�'��F(��-��.C�e�>�77��v3�ylG/])��M�
���y�)/�cb��4}��=�����u�?�IF��Ƴ\c$�R
���k`[���^��U��d�A��4<͔ ������x�iWjt�Ƥ�QHڜh���-ͺ�$â��A�	.���Y�58DHu���p+��0��n���ґp�?�����p�ȥ�D����Y@v��z�0��������s�* �2:��;0����E���լG��`�K����͢��gB2�L�<�mG��|�P �����>:X@;�J&Q�40f����-�o���Ͻ�F}&���w֕K�'���'��Q���R�V��	j4X�
���#,q��U���`"2��z]i��g�߅�Oe'Q���
�0!Q|3ڐ����s��Ȓ��`j+�S�\��i��X2�vE)z��ν1�4��!���d|�[�qs��i���My�@j����g��XD��������o����� �#>% >�z�X�PI��g��@��N_/������y���%
�Iˠ;�w��z��2I����<�A�̝SZ+�pi/��~Hם��>�w���)ԃ��Xx����"�iƗ����@;Q�,���+D�L۟��2j���$g�����;2�Z(���=$�e��͌�Tf��+�ɚdG0e��Rl;���@����3)���A����b�ɪ�r"��&�X�`@z�x�iLwLa�,�K�1m��mq���g����r��UvKi¾<��rv=��B~`��3��1�������Ș���fS����B64�Z+wQ]�|�ngM�)2%qie�wh�8�C_��=��F�8i;��t�\5݈�[401���׼���t.�ʀ~�1�z���LHdW{����Fފ�Y��F����>����n�aT$Pu���
�7#Y� �������
��J5��Ry��N�- ���ڟ�}2���y�5�A/�H-��N�TZr���{B����[����o��Mb����J� �rn��D���#�2�v�;�ǉ�����.�H���s�*��ޘb'H|,m@�VKo�vW�\�Ȓ�)C�o���1�����Xڅ���EQ��'p�T�!j�Z<��Ui�r�D(��ת�ѝsg���5D�����l��B���R'�����m�a=�� �6j׹�v� ���,�3�''�<��,> ��n���2$��w��"]x��n�����M����>?��������hZ���6@հ�2�_��Tj�p���e����$�[!�-\��Q�,E#��Y��cشA��V����F o奛�Q��5 ̔�D��!l�t�W��
 �UD�}F?�]�[��z��V���G< ��P�LB0�,6 V�f�"伟َ��,Q��Yĝ�>����4�<�L������CE�(4�^��_��,�|�&Tlw�Ɩ���ő^�\w�"ӞX��{iC��7��w�v�V~3[8S����m�����bW>����E.8҈�7�V-A��c�Ro�%R#��$�;|2�\��6D�T��tRhӸ�)Z��=�����7�8l��B_-��0Ս�}��v��w���4���D�>.�^�.�e���tǴ�鈫�Tjhrl$�̖)-�t�o$N �	K������9�	a��g!��K������v��Rn+��	R��S���1�E�N�i��>�0��`6H}ca����e,O�i��6z�>�H"YP��e0�G����d���xH�Y��i7nmT���i�9R��Z���v(@;Śy�h��Cr��)�u��G�m(�����;���iec��l�:��uVԡ������a26�r���F�^8�h�7�Kkp%+!(_�=�+��݀�@E��eh���mS�$��	9K|sz�x�� 0��C<G�Q8]�6(��'L~�K�� ����JS�jp8Z9{�v��ߣV��(`�� F/��#�$'~B)��t�u$4K��	�uK���d��� �o�x8[*�P+����0pU��	���vV�I� �2�� �	�vW�e]�y��W��`���K����ٓS�G��pv~�Bi��m&�n����!N�b?<��ިOw�$��l��:+;b�κw���ؒ@���~d����1�^��Mښ�-Lr{z����N��@���m�G�Ow-`���z/*���~�'��JM���� �;V*�s�Wy���#Ӳ���S��qm��^�t6-��Y�Ė�/q�"lN�U��u�_�f�{[����ؾ�$�F#"ղ�]���*�/z��vź�1y6�3@[D���N��!�i<�����������1kّ�G�Dd/���e��BŮ:�*fsg�M���q�c��ǿ�Xu\���n{�q���a��$�}�7
[�ҟ(m2��4��&\�O���y�䝰�0��jŵ�Έ�װ���Cj�_a��>Q	纓.��%z��I&y��p��V�R�Z�\ߓ!mS\���<Ad��v�e粵b&�#Z�j�	+W�'�c��RbF��c�G�q��#�"bs��N+uJ�l��C)��\��t����|ǮH�do��ஓ`t$
�K4&�n%�_��8�K���AlHD� PG�9d���z^bԐ&��,����Vɚ11%dH]��˯��`�����"??F���x��&*E���=���
y ����۽5�V�I	B�qf�t2ϐ9���D}e;ߣ��d�sIP�T�ٕ���e���C&}��g*�Qt��H������G��Vx���_�:� �����A�k��BY��=��"��Ŭy��Z��˕��󟤇sl�%#"[d'�k����6��J��NO:���{໇��^�K��+�����#Iܥ��%��Nmy�I���I�bs�:P���MC��G`�«��ٶ����.�N �;R��a��
���n~9�x��^�.�Μ�]k���B���P��3�.�
8��j��Я�2;A�d�6$��JZ�#�6�|)�x[2O�I0�>҃�b�i#�L=���i�Dt�����u�mM/�Q��]}�en�q���(��� ���X�f�s�K�����+އU�Q���v���@��L�􏢺;6�D1�sQl��;SD��=5��$�Ow�&�����X�m0�ɓ3V�g���1�}~I`���:��θ�W�?zŕ��2�W�G8��ޢ����U>�A�̣���1J��#��
�M���C�d���` �k� B|�M�2�RA�*aýodO��k���&��v�ճq4��y��+��;�t���׹�A��� ���"@�\	�7� �q\̞[l���c�8�H<d��ֈ<7���PͨH�e���iRkꜭ�N(tAhj%�$y��c�I�/5��3�"#�.��������  �e���$�|Y�ȱ� 4�v;�ӝ���EoK����:cY܃MPRgM�W�Z,�_C�� {�f�yt�I�������mƬ�)Rmr��j�#Ɔ�����|\��j�k�]W��oϹۘ��\S,ҊLIǧY��Q�.h:�$�p�4eU2��+l�\���f���wG��T��Ř��I2x���B�����(������yx�&e	���W�F�6�1[��Õ����xHb=�+V.{�/�����UJ�^?���۱�^ډ�1^~^]o���[1���|���	$����"�P�#%���[��W!m�����˕BAaښ'�X�;��L2zk�J=&��R>~���O\�B���A�tӈ&Ɣ�2�'���A+/��5lgh56�~�EF��	&�2=_i���$S��n��-�NQ��BXBڗrߡF�-����>�����هVN�{��0��w�ߐ�BRf�j�[߾1gE5tH��C��v���c���r�ƗO�?M�P�������� �+|Md\�����5n�ҕ2.g)Ԣ��]��v6� �%b�$(r�2����m�'[��m�;�C_~.T�\�`2u����8�K;�}��.m��b.I�u(�0݉�����LBzS���&&�˸�����@;��3K��3�F$d����j�*�΍�e. ��\Z��9S�m�c�K;�՞3�̜���;A�mZ���-^F��[II��YYwR��wǒP_Bqw�_ߌˎ����k��� `�qOc�B��YY0O���@��t�o������� �
 ��p�*�1���5�ɵ<�\���@���ku@fב2���b�艟>'�ǽn=��C�u*B���¡C�����iX8/�C��>�h�>��g2�e����0!��2���<K�C�� uK=î*���N �%ثm��u��r���~��,����ʒ�r�_�8uG�j6QG�7�y~�0w6��o��	���m�v���� �-�$RDj8o�_DG����� Wl�jP2���|x��E���Tj��r'�#AF\��CI!�ju��Ca/�e���o���qa��v��Z�.@
c�j�9���h<��QP��Ru3M[n���J+7�t��/Lk�[�����#0u ۆ�Py�AX�2a�蚠��$�]CaDY���,��mA ��*�%�4��2��^����n#O��\���E1B���9�*[���
�l�64��^�E�Q��k�}w��� R�뱘��0�f!�86����3Nٸ3E�[��P���7���l���g��o�<��@�֜쑵ԅ��G�οFN�����{t�)�a���_��C�w���F��|�~����z��e@�շ?�z�z�Ө��%J}�\f�2<�!,c7������6C����$�����������0D���R�`�
�����tZ��I�#c��X�܀n�0^$˶��+�§�ρ����SE����R!	��uD<r9ןP�ѽw��$�vU3h'h�l:���0����2�S�!*;M�K�6#�7�����$�l�W���.��0�rÕ��Fލ!SP�JT���U�fĒ{@�����q�L�pR�Jh��W�C�|�{��{r���A-v�#+zVB3�nS�Vt�����j}8�a���ݢ��� k��t�]��։^#tĉ  0Tג��!)�G,���\�|�@��i���ցߚ;�uL��D�C�J�L�A��Tk����mO�>�	ɈO�3�'y<�~|l}��ؚh�r�l�ZS∙���	k?/i�� a���6�a=ȃ	�*�Vj�ZV���8�ՈL������D�& ��P%����%x�$��@������2'4��m��5��u���HA.Rf�ߠ�)LF�ts ~awߢ�r�x�1�v�o>3��$��V.�s&�O��OL0�&wH(e��Q���e�,��Y�C��
\���,`��ʲ���<��"<<}���K���n����C��G���@�~�"(���"Ԟ�=�s��/�W�Lͫot��x����!to�LsdtV����ݥ��_Ħ׫�P}?��&-%�=X����-|;�+�'�������ɯS}�8*P��2QIh�5���Ы��,e@��+j_8�B�k�|V� p �T��c��HF+9a-�g%J�
����_����+�������9~�ף�|��*�ўg������K����qtU0`v��\'{�D�#Fu��DP8�)CB2�G��+	l�`z:ׁP��A1A�;g�$}�Ul����BW��)��j��1��T"������*�3o�^�$�>��>�v7ܶC��5z��M�����>�٬kJ)ICAvf�<��|T�cE�'����	xB�r��Ж���e��oL/_/�����M�������_s)�.&Ԩ�xh�[�b6�:�,���Sy��x�&�}�o�Vb�k�9�]�K����f㩥�����k�KV
k��_&!y�b"�!W�WE�/��փ�����óE�ՙ[܈X�|_s�6�rq���"�|�{N�r�˽�Z�"и�;� �NO6!�'~��j�Ͻ�?�AZ���U����wn�4Xm`���2F���F�%���k�*�͟��*�m�(�t�Q�;��Bӽ�tI��оe�,m����>'�8c�KO�	���ܤlZ�|�>�3PP�Vm�J	uL�Ǭ�7��@TMވ���sa�<8�
�须�Vsz�z3���V�\7q1��ޕAV���&r�.z�]vCY;(@k�1��M�heLY���T��o�?���@D�D�im/����rj�hR��'��t�b%�i����{��d�d|j�NdKjT"Hʠh�b�S��sR���;H�U[t�~51m�Ɋ��_���=�l���0�:uł2���QU'I�%
��+��i��0(�]ズ[d:�.���4Xgm�?����4���������o�c:�hࣤЙB�&�#{�V�"�<_Q�8���ٍ�K\��H��K���k��ɂ7��ޝ����[]M7�5��s��z	�I�󓘾�(�چ����.f���@�Pb���%�S���a XP����õ��o�^ku���騃-����\Iľ���p7[�� ���w� ���j�.���G�u�"t��K�m�DZ�V��\8�r��)�HW��sJq맡�2O`l���7N�8� E)ڿ(�U�l�q�is[vC�����F����M���&�!��d����1��{Q#I=ug���85Ti0I�#G�|;����'�� Ik?�B6�R�
j8,�jR�a �꠆2�&	Ԑ��;��}gp���>�_��Dlc���/lr-D����}6�IY\�$ =��w8��pR�����`��d�\����]��B*�S@�U��=�mv��ܞ���LH��%]nZ�V�?L*'Gl/�!��e�[��TH�I��mé���#� ق_���+��%Z��R�����E��ƉFg���-�������2;�u�<8K���iiQ7�L��D�grɈ�k� ��R��GdM���+���
�y�j�s���@���H�����������0&]��K9����8���^[\�n-M`ҥM��,�ύu��^;���
���w&��ՙ�9G����aS�Oj�x�:�<�Q�׵��P[+}i�]"Y�_�Ê��/�Z���uF�%Z[��Ś������}���ϩ'=�_{���KQ2��k�za���y���\���&*@���l��\��U���=[�7���彮:w0{1(��e��� h�%�@�L�'wJq���2ޔ�S3���Z�)����5��&C3�B�n�nV��c[�H�@5��z$�9L��
x�9��ú�=5���75zCB�N��:Ȩ�)����-z=�+�Ƚ5���3�>J�WR��QU��m���M1J&7	�`C�q�#�]�$�ӷ�Ԭ��z�qg�g�3�iä��b � !m��Iwf�Y
���ؐ
�n�ӥ~���ً@�/��:����0$�u� c������Xx�#�oR�K)�"�kH����k�Q��ϾY�����P�>��ގ�8�a�_l2�! ���9(�_�m���a���ќf�6E1��ϊ'�sZ��0!���g�[~�.��%M	����� ʔW�X&��v�_��;�4��n��zN�Jь,l���'Vz�nkn ����~�W���n�ސ]���DJ�3��W��i`���-��k/ф�gڣ����@?�ٛ>�ܒ&$V��]��9���6���L\ IְOT#~���h���i���Ȯ���� �ϐ�'��U�
:C�	4:U���^)�~m�M>�Sf���Z��|v��ZG�%JD���Qp�6�������L��kk׊m�lŽ��I�"�]$h��Ĥs ƻ�fe6ݵj�X�t�JW�-�Y`MS۲�C^�w�Ǵâ꛽$�?�>;�"�k-_����u����B�C��ku`~�%u~�{��V���xY"�`��V6�.J5��@vu�\/H,�9��"���CDr&��>�y�뗠qE_��,)�H/̛��ꕛՍ�b(Ѣ�ޫ�0N6����p)n�(�����z��<:b�~%�@����U�J���Q�.DG�^��ڜT������5�RA�oq�}ת�Y>�ɡ�P�6�{�������������;%��x��jn����Ģ�pYg��2�^�cڸ\{����_�H�{b�%H�u���"O$_(|=wX_�Bʟϻg��u�N�����
������#��>�M@�ޟá��
@}�kw��m����J�P �?�:B�������X5/����C�4�N�o�n2hԪ�(9J4�a�6��QY�𜕼ZuY��]��*%@��F1�t�����6<R���p����pֆ+Y��8�Ϥ@����JE]�����|��-p�}g��|�ѻ�if����z. �z�qˊ�)�ASډ�V70�V�AN\���ˑ$��c�.��&��wE�5,GG�p�ɆΓs5�k$�U���(��UlLM,��X��m�lW�,��B�1�[���ZK����O�����C� w���m(��	��$��&���gȷ�������U<�M��aPd��®�����Ꮪ+:��_̢��vW+��{R���,Ӫ�H}�+#c���,�Tq94�~1l�����S�gu ��)�|���^��ǘ�+@�bB��5�hϝ�.��K\�:[e��|��(l��r�W����/���1׳�s޳�|�ۆi��)�,}����Ik���`�����D���ZI��@ek��&�B�����;��<\����Vܖd�e�St��c;i�d榚�5W�E��Z��' �HdA��ϓ#3�!�]��z@+x5��祹r��-Tn@�ZY�O�X����Q�+e��e��`֗�!�él��a�7#i"Da�qq��H+�d �x�g�~g@MF�j\�]��m�8�T��(;�����VH"4���	�/X�ە3��د�]���(F��߸=�@�Ӯ��M�����MfS������	�2'��ߌ�sN3y|�3#T������}辣b�.mI�O�����$Ѽ�!+Jv<��n6m�/�����Q1p�r�)�s"�7q�TAX.N����B&��X�P�D� ����+���0�gO��E] ��xN��L��К�� �����0�V%x��(���@��6���9�|�X�Y�eh��1��#$��^��ڊ��8Ԟ�y�S�~���iAOZ�]s)�k���b_��-$L6u�H׆���j�b��mI�c�21,8��ǩ8�+��c"' �=[���d�5��X;�@0<��*�ӂ�a�^9-$q�.'�HS0��3�U���j<̆��fa��:r?6��dP.-�`���rż'޿�X��7OK�P1
 �ҍ��O]���M����;M�f!���,�x�c�Ir�N�D��BMQ+� ȇ���~��
4��Þ��s���^��(��Cg����H�Y�΢��y�������1�)\�J�K��{�0f�C��ɝ�]��S��L���h�k�5��m�'���h����N^l$��s��/"�v�����GU�7!�Z��"�ID~V
=33u)�N�z���c�n���
����OZ�6�\�w�W/����t�猉zh&G�3i�b��|��
�*鶝&U�5)�*�D�I����T�6��b'��fї��a�4���A�����D�S��LM4r�0*��t�6"M�@�g�Dg���/���n�����5S}o׍P<>�A1Q1�A̰�ֶ���;��KK�5�`�
���Ձp�R��r�1s\������r�ര�[�GLiI����!�\��]���]����2����+�.�	���[?�&�^�<�$�*�8�YU6�M��������5��p��W��6bPc��wB�򎷿,%��7���t��2ʉG��R���)g;�p��M����+�*F����Ni�Qf�%f���&�ېY�����\ژq�Z�_�C�}���0��~2,�tv��t�.jZH�S�6��X�OL��X2�u�ܯ�%�YC�c��Bes��oP	7'�B�W"(o�~��h	O�UR���[�����>���.�I�G�>{�R��p��%fY���]+uA8$n�$:̝s��yJ6�+�ʲ�{-@��i��hI1��32U�Gl}8X�@b)���v��v�bѪ0t�
'W�<�O3 �2)�O���׿!Ԝ��Б�����5fI��!�+��C0-�"{�k i��=�!����,��	3��Z�����;:ҋ�b.#�`��0Z�V�lk��v�!^�ω��S���Ur���C�q�����xnW5�?jZ^����F1!�Nh[?cq,6�g�?9����`��X�E�;�����6�(��H)X~�����X� �`R�I�t������ߨ��-�����ע��i�k�[ئ?a���/GJn��c�(���ٸ�mQ�dW��,4)���1'�F�o����ǧ�$�7,9�$��Ftv��!/� �v5(��UȘ��XD� h=p6rWa�L�#��6~�:�%���~�JZ��7����/�.�&���������4�C�^��&�v�5.��Mԛ���$�l~b�QtA�Hs��,J�Z�=��N5��J�9��'H�Z�ada�2m(���,�OY�i��<)��_V�FLK�����n����YI,yt����_������.�Eg������˱4_�у�λ��f�+�cF�iq_s@u�޲�4B �=3i'�w��.(��7s��(�Y��<f��W�d��9�8e��p-�*�2aҠ	�/j�[ �SUR�#�3:���2��+��Y�����\�0F��'�H�l$�,�ɍ��j02�x\�r�: �������	ع����.�z>�r��<�Q&4ϞB�����2$HU��BC[ �Y��3�/�(�E*�]�S���#x��yIG�gc����ϓ�@r}eD�IE�k`� X�=(�j�t[�%��gd�d��d��p%�ͻո~��U7�s�z��&b$I�x1��\�X���`��)nQE�����$�hW�_E�v��ƍ��}�c�p���*=$�p��h���5I9�-�aiJ�dJ]]ɼM\��	2��u�s&��Bv�tB�nr����sz0>��T\�ҼC<w��!f�zcp Mon�QX��ʽj#+�K��
7��� '� �3��M( L.c>�k��*�Q+�u�P�Ϻ"iH�s쩖��L�g?��F��"�cQNHފ*C�|С��@Է�Tp%V���	-��?~�e�r��:�H_慵se�:��&6�3*>���ň#�(���
s�}�8�X�����8���$�)A���o�Ez�Ȟ.�3"|.Ά���F|�VGp�A��Mx�W� ��x��ن�?؞e_V��8J�	Ia�W�W��NG�#N˕�s����-��Q���g	�ɘ���5*?)iy��-9�H!t�3<��ȃ�Y7�$�!�Ypw��ץc~ޜXHN��O���#��V�3ռ&R��\�i���*�#�+/2v�#�
u�NO7��[4�傼����� �a�%�C�q��5�ݫ��b��lD`�oHYX&��QpI�ʘ��UD��TI����Q2fs�p+y����vԨX���A��/:��~r�w��,z���a�D���_d�	��B��#��$���;��w����x���ʃ�
(�d����yq��Gkgo���;?"���G�hY3�e���BI�������3d��A��r����^~��b�Z�c�@�I���ق�w��6wEz;�q-��H%�M��`�[�����W����4����������������S�����1A3/-C��paf�3�x��M܉��ҥ>��S;�+V�71�J w-5�W��C��O��f�u���r�e�0��Ha$����/k�K���+�\���5��Z?�#�g���f��qr��Y��]K��c�G�J[�����)>ӓ�&"ٳE�C�o� S3)oaV�<�u�_,G�ܲtEuXYZ�����:CY	�(����Lz��(��o��<��&����g�Ps'�H�kL��S�uR���C��ׁsډޢ����+����0OpN/�m�ֽ��ы�9�t�(A����d$�?k`�	���
B�U?| T=��	k�;]�U����3��Pl��c���P;.Xc�L�4���`��S!vKom�C͏[<{���L�̨���ʥ��Z^���Q��2�4�ܕO~큛�&�.�e_���d:��p@<����S.�#6#g��v2��{�i�_��۷Z�`:��6^4<��rL���
����,�Ya��(�o�fk���tD�!�s�����ǂ.�t'���n�C=���1�K�������R�9��|��C��l��X�ԞEA� �K�\]
z@���q0�s�2�ȝ;��,@T�<EpZ7%0�)p���m#�v�6S���vwqKnq(Ns���{��6uI5��V��&�z�,����6?�? ����k;$%����l���uu�ϱ�~n�HDeo������_@Y��Hʔ�`����=�l��P7�,,����\���B���2Ϯ��vfi=6A)ĵ���nz�<�-T겠���t��փ�-��U'�T v�[HM�F4"�\��?�&X^�"6��A�`ȶ����#�fɜ���M ��0.<Cǧ��!���L���jMa��:���9�U��O�����XFSGJ��}xiT�S�~��S��5%{҂(�N���f+����|k�&�6ܧ�����E/��V�gE�c_y�ﵤ6Mr���8n�n�Q4��n�͜J�k�B�F����z~�����Mc�e�������{�\�>��}!�>R3l�uYmFȺ�/~E��p���>>6�_o�����]�w'��7yi������4M�n��)V�8���$�_6u�fb�oL=`x�g-ҭ'8��?�d#"��!�"�{A*��g���9[���Q9/�f��"��`�-�wS%�/�an�wL
��a��Gm�7�*	xAI��x&���_�eb�����j7��sE7�@��.������9�~����\�>xj�Z�ⶈ
� @k����G����X��K�n��EU����@M������u��	��	=�� :�� ��W��D�F �a��v�f��(hO�������Gʸ�}���Bǖ|HU��|!���»��7�?���(Ձ����%�_�3�|{���,��Hl1抒���4�B���"�����á^R����LC/g�4uF'���*���{nK�0)����qs!h��i9Z�F� ]��`�����~�{��q>J���:5�"���1��/k>��m9�? t�fCc��β�oȵ
��9���Y*H�0��[�>;� �d��3b�����,�Y|���3��W$�c%I��6:�~�J��O��g?�y�����!�;9b/C���:��U*K��m�#S���9*�9c'V(a�;2	����1���<ݾD"��26�lj� ��'��bNuM�5
,��N�c��r�r� =�W�ZKj�	��v]�GJ���<Œ�K�Q��]��7�8yUL��q�_|o|�g}Z;�TF�ȼ!����<�����G4e���d��-�g�M;(Yx1� �'���ʹ��D�K�� ���[�M҆��a���ky�h�x�2e�.[�V��)O�"�21D�A�;r���Y�L�cE7���M4����;w�{�s��
�)���Mi��,���͡�C�6��
�>�~��<r@��\�k?J�iL�Cn��]��w���H�ʽ0��>���#=\�6I�ޒ�y�mK?�!���$�>�
&���5�q��Z��^�2����Q����uظAc�I	$�A��$&$O,�8.����^�t�u[ w���7�CƳB��s0�NIal s9�����mM�o���h�f��W�^�Mh>��"�9�T�'��Ou�tc�$+�����?��Yd��� ��tʳ�<�@T��L���8ߢF�8ڹ��[���W���ͯ@1W�b�jb�����( �F@o�4%kd�T��@�j%�i^�f��n�j[�&������>�F��\Ċ�ܖ�$��-��+�Vȵ�!c�k�E���v�)q���S	�z�M�`����D�z��npDB��NMy0�;��g���?>9ӣf�7����y�->��a�}u�� g�-����'��c�4ׇ.�3/��@��
0�X.z�n�+����K�*Mc��0fO#j�-��v`����mn�5Tp; 
_�}e]M�	W�?��dH���e���7��S
*?d��Ι7L��ߕ��$�V�R�x&��u��Ve{��n'K��)�\��n���4�"��a����u���jP��oFh��X/��xj�.J y�w�
�H:��C^J^��s&�K�e���(ޘ�>�+���2#�b��6��8�\ض���,�	��!�����ͪ��!d��2�ׯ���{]{�g�	 >8ȋRpv��U��#5d�=gi˧��X����j��!��i���ݯ�h7�����"敠���Z$��C�[$���f|���-.��Xxaz�VMcr�hD~�a�2���ַ���=R�r/�6#g���W����dꚸZ�$ʔ��`���0���x���h�YGv�{�2�������_y�i��ⲅ)i(��#D�T&�Tҋ�̧�`�q�R�ï�%����2�7�$@~���`o���J�d�R�>���!<otҹ�k�^*�M�eԫ�%6cw���[<_&�bb�'es���YM{��b��ߺ��)�:�gY2=h5�峿c�a�{OtU��צ �t�G�gnn�w$ֲ���3N��0�C�TZ��w��(
�J�Ҿߠ��.��6E!�E]v�9�L�gB��dVAT�ٕ�pBy
ǣ���T�tӟ�H�����ɠ�8����1#ؒ}�����w+o.����8?��?�놫"t!G1'u�j�l��jW��{t&jo�:X��w����`�TB�*y���6�5:
�W�\		w�dh�����D��֭h����L�ټ<�y\@��x�����2
ć���;�>3���(e�a��l�/�����ld�I��P��fH�*����x~��O,в��׸���^h��O�b �Rd+e �L���N�;I����cUΈ=RFY��T6���ɿE��Z��z�!�VyV;F��)~�!U�îY�)���.�
,�qa�ʯ��[��C����Zsh�� 
FH"t�q���w�p�"�������G6�^��&H��g�-�����Z'c�3�.7���̉i��M쭺��J��e�T���Tn�S�Ѡ�����r�<+D�J����.��%��܄����$MN1T���W��������K�Gq�a� '�0gz��A%X�4<=�uq��A�o�U������G}YT�e?�.��e_K���[-���v8�+@P]�zB:��#6�y��t����?�3�@�:��0J���b��e��f� w���jե��J�Ny8����D~�ZLb�������GG���7t�S��h�̯τ��#�cl�O&���յ���H�!򮙹
�c��g?��X[*����}DP��{?�п&8A��_Y�':D���2l��j��N�Q'0����0B5��˒�H��
���&������3C>��'�nV�0���F���zR�&A���n���z9��������F��
kl��u�Z��W�J%������tYs����M�7��"Ԗߚ���+ؕ9ܫ��M�V�҉Nz��w9{����ʤ�K�®}E��"��vu�c�F��vu��3<��yX������7<��H������� `g�1	�H�.�!B�{d����2r��h2��� ���]Q}JS��6?�h�o9~��;����C��["�qj�+�L�u�a��Cv���sL���g71�l��U�e@�C(���]bC�..b����i{�i	 o&'5��H�\�m�c��O߻� F@r�����؏#�b�L����8M��NY����o�p�W�����u��ŅB�`�L��&X��$F���ߟ����+�s��&n��l)P���MVN}@��f�}5e�����*�CI:�U B	U���K��<d�_0K;!�\���O�0G���c�����_B���]���|��䥁DwX,*o���lį��T�pIP�,�����yA�����F*=݌ҟ&�������֘aR�C��!��In	MW'T�ǮS�2�w�Hl�����O/���a@D��Q�MrjR!������}�M*�a���]���Ad��W'� �ܧ�t"5�+����F�b	�$۾��.�`#����QMk��-
�xiG��4��S�ͣ;"�c3��cD���1��Z: g�i�*Vz?w��}��J�}"z�:	��=*��)K�,�sX�Dk�Y��2���� ���ä��`C���o��u���zє�n�j�]3?�\�.'j�82��]����1�E�/�[�����3Z�RW���+��N#jm�N;/������� X��}+в��-{������K�!eM����ӯ�Y���kiNU�� Ig��cR�$�� ��}����ߴ�L�>	�VD����LY5�ڵ�O�q��[j�Y���$����У��(N)l:�����D�m����!��_ƈ)���Ȑ�u��3���߿�%|v��d*i����e�1o#�!�$4�|���֮�C�o�JmM&W<� J��L�#�R$9
���$�ʐf_�h#Ӎ¥`j���k {Ȥ��z�إ�&�Je?�d�R�'��{�ƫCQG	 �z�f��$���Xd��C����O��{C���،�[f��x(@��D�$��M6�W��J�<��E"D��L�����̛h���d{7?�����O9�F��-�2�:���ኔ�Yy�c/!$����JR���(P\�4�����ﴛb�_�q���7�_��n�] %���s���i�-��b�S�M0%m��;\3b�}�X�~�B�?8\>K2Ѳ�s%okY�$�H��4+p�qƔ߬��!�Ί�}l��y�U_I�?K�汛��m���Í�@)
Oo<��OK���d��SӀ�\)^��u�D`�����!����k?ԭ=��	b6��%�q�HC��V�lh�� CY��B<M���$D��c♱&�Sk��>n��7�t�d౛k����%�s�3KJ�OIW5t��2��s|���b�J0����M��W*��uh$e�酾̭�,��y'<on�ޞ+}��+ʄ�V1(��l.��w���JћG�sp33�ԧ����u����G���n�mZ���){J6����]�_��H�H�%�Q2������ꪩ�[M���*�(�ݶ��Q�#���墱c��^Y!_J���9ޒM�E�,�D{��?0Dj9y�*��bI���q�w"2(I tA�2��P�d�=�c=,��vQ���0� <�[x�g2���Ƈ�\��R1�YS�ۼ(N��GP�Ѐ�C�7�T �o��~���yc,<��ʠ� ܽ�֛���ω'm�7k�)���rDcрV>Y�N�<�����TγSO�~O?雅h�cVy-��%��B��,؈�D֯&`HQ9r|c�(���iX���r�pR��í֣�.NNp2D鼤�h<�ř{D@	b��r�����k��x/�x�U���%ӊ��@`��'*?n����n� ���فl��U@�n�B���l�a���93�_���Ar�>$��ն��@�N��K�	y���@�+���L�����=֣ۥ\�؏?ʯ!u�J6��CZ��OK¦e��-�5Q��84�LMta`?2IgVbiِ���&�� Koz��J�;MG`ɳ�	|��\>8�UJ��}���WV?�Y(�+v�ϒӰ3�.mߣ5�k<A)\�I4�}	1��m:�9��X��|v�\�g3�����`m@�T�ƭ�2�R���GZ}�J�97g� {��o���3*QrBCa2���*��!W�$(�~��}�^c�J�MJ�]�Gwr�6�������,M$?���R%�+��S���g�Y�����D�S�v���,�v���i#��������0�s�1tB�Tc��9S��<��ѥA�K%�Ƶ��J�0���o�χ�덑r�VH�+�o��e��YxP�V!��g�֓{��n��	g��Z�0����@>�V���nzE�[Lϴ��b�7�%�9�R����o�kOho�����"�p��22)�����'�����e�8D�j4_,�!ON����I]mG�ĤNt5f��r�C���J����,�O§��l��n-��$��fo}i�R!<J�C�$��>�h�>����h(�T�(��$����X_�I�3�Y��m��k�<��Ŀ�����R���T�R$�HR�I���(f���/vL� �����U�(����3-�a:X�u�O�$]���D#\/ɽk'��K��"���e�҉����u���0*�A|1I�0��|���ճ��o�J����!�n��V5�Gӑ���dB�2��*Њ�x<�,-8ȬM��$��T^W�;k%꒙�I�q-��v)8F/ ��I���T���"P �_'+xuՔ�
�S�{zIu&��-�k�5�q�rBj=� �/h9�����0���}�A/V��J����Ql�Q����� ���d7�=ݾ<�b[d�"��vgM�PW��k��L��Ɗ#E���wB��b77"�$����a�GhI.^�75����4��|�v_������/*����DA ^�2�Ϩ���U�������ɘ�\d��	��C�R6J4u�y����.���ZX��G��Q/M1BpH)�<�L�;��x�j�]u6#V�h9_���bTS���rAL�����F;7�SJ������9���G�@�	e��z��iF
�b�D�^�]i�؋_��k��Y�j$��ܱM�0��;�?�`:1p��5cO����L����aCTV�e��L[��9�Z���2+U��%�'���>��������#k���B��#�g#]��l��T�e�vr������k�ާj�����2 4Q�y>^7oj>ߣ�׈���Q�D'6���Eh[C!�O�25�enV>�lS�I�gE~�*���'�;����AQ��#�u꟡�{c0�C���,2���C�D	���0<��q�&�W6P����p�-�E�&J���ϵy �s��W�-�MC��'%F�-�H�fV��"����z��r���ADF��Q�[]L�}N*�|��R��.�&����d��K�`"=�}�w��:��欷(�&�����׻s$^��� ]g�%�i���)�x~��~��5	�r���ejk?��g�GPA{Ѵ;���+���Y�(�z��Hֵ�!]f͂P�6"X��uR�|{e�Gq�5�¼�c,8���nڤ.��
)� ����g�H6��ϫ����59����u�~E�;�"|�}ͽ���;~�p��M@��%�17PH�����	ԴuL&�=��Z�Sq�Jno^!�m	fIL=���F�.���A8��s����������X�oF��4(��(u$Uc>�;a�=2 ��:�c�*^�WKl�;A��>�`2�Q�.� �"%�R"�aJ��
6���+�(�$c#���]�A�"ݒ�d�~�����Sjޚ�.xx�6O.ޕ�C-����<�����1��m���K6[1���ׇ�F4��/ aeP}�:���了=��=���n ;���Ж�:���6�U9���y��t6��|3W��^�1,"�=���"a7��I�(M�z�1��?:��Z͊�,���A�݆t3`iN�Ce��璢 !M�Jv��Un�R�x��$��ĵK2�i� �$�<���P�&�
11�M���2��|D����>��a�P'���3�x�r�C|�[uU�FW��Vf��LkX-�C��Aa�G�+׽|��ǨR2qX�i��\�#/�E{�R����Q?�[�QL��b5��dKO��	��:���&	�v����+b96����얁Y���A�����s�+��Т���l~H�C�����cd&��D���XGP����L+�!��޹y���!]KU=�*h�n��0 2o�����X�o�q�h<|��@�\A��|���'�#����j�[WwaJ)XZB ����'����*�zi���)8|�&�Yʫu�[����l#ޚh���|1m_>���2��.��8��x5t�y��܃1�Wh@n蕦C������X�nT��L[� ���p^�7	��]�'
�q*^׍�iSɜ:�	����o�J�BLA�x@��Lg���-",^��U\I�V>.n���<]D�A�i�Z����f�}�AYo��)[A�;N���hJ�~o('���X��p��R���se	�$�=J$.쭗͎7#qƣl�8-� f�7B��\!��%64��#H"-���]q����r>�����V)��F4+�h�H�X�U���Wb.�r�`Bt|$�:��p��]�iz�'q�_��ջc���U�!��׹瘀�]������i{?��X+8�1�Ld��|:�c�=���@�T��L	4v��`c���M��FZ��5�\��#'ɵ���]���34����R˿�C�*�#i��,h8��ۡ�7pi:"��َ\ �����ՇeR�!��9��O���$=����i�����َ���(M�<;�����d���]�D�&Z%d+6T������t��t�'�w�z|���t��H`�N�`!�;��^ɋ�*H!:���i�~�/��k�O�9����F����ʸ��v�����q��y{&6ɉ�տ���\�ˍ��z�4��c"���n��-��K�vSe��K�)�f��]�����K�8HgO5�Ͽ�7���F��(�L��hU���%��"Zd�'*�'�Uyܓ���e_�[!S7�n�y�e��<Gio�zV�ofF��u�y�{���ąU<w��p���;9F��/;R��<Te%y������Jh��o�@.�{�Qh�.8�����(s�/"����x����'�xiZ=����M��#$ڒ͜�DM߉)�\I��ȅ��p,v{~P$��cǈB�������� >7\"���� S�3.��~���=q �@�4$A��MB���>�u�e�����'��5w93�P���2wa
T�ktWp�Ф�m�@_�`���Ψ託/KTY�s���_Q�/���$�+>��i8�&�����%!eܿ���!��3�=�DYr�zW3O����>�&��.��?2d-y\'3��E6���S�vh#G��?�S� ����2p]�|�FIT�٥���z����c�뛀٥��i"���/��	}�O���ʣ6 I7��ǀK)Ƈ����La���� ���`Ҝ�V�a]O�H���Ҷ�C5���c�vM�A��;m*aJ��^��X�􆚎��o&xݻ����uWlf��ך^S�0+�����?��*��642-�Dڍ�|Ze��v?H�3D�+w�B�=0�"FqC3�� ����G����w���g�`�,���TKH�g�J�7}qw8sAj\^c���7����I��ڤj��";�D�����1i��;"��{�s��D##���!�d��C�E�a,rG2Fx���a���Rgb�nV���\�d����I��ٻ Փ�.����PƤ�Ǵо�6�G?�m�����?�-��g��hی'�#�/Y����;i���&S��*D=�S�`3S���)#@�C@��j��]�}��ޥ�͒z\|�=͞���
'�W��Z�Ș�KY"�߉��Y�E
�i������W�����=D�\��( o4_?�i��@�u�#����~��Z�^�6�	�`5�;��O'G�#$ʭ�7�A�G>�Z�#EE�Db����l�H��H���	N���b���_���}_O�-
������
IS���m�UZ�@)����;�G$�Ï����×�ʽ�̂��6:��S�R��D��ɳƷƶ����d*]�7DO�ɋ6~�]b�}w]�k��2�T:jL��8�	:�ު���V�p��
���(%��ɔ�HͶҦ�ر!������O�C>|ݯs�(��l"85 s���OK�(���8ؘ3�~���Ql��2���}����#�<�u� '�m� ���r,�1�h�xK��&�?��iUU�b�����?�8�e.�r��3�=�n�Zǃ�$���ǌ�
�8b<�0ʾ��6T�մ�'�:�,��$^5)�S�F�E
��}(����A�)�exj�y��Q�C��q�|�̜������bC,�=1���9c��S�G��#����y-S  ?�# ���B��2\/ߍ����`���2�|WۢPp���V��#aҘ��]w�_�F��d�$|���&�k��9�H~����k��Ei�H��CW��]��cr���]ˎ|�����_G�z�՞"�E/д��+b|�}�@�d;��F���;�AQ��r@f8ي�5͎�^����GG���p9��瓡?@�K�k���&h��Y쫳U�q
󲊎���l3�<%�����j_�&��"�=Ɏ�����7���)�+�c�(���g.��Z_��$����� �0�zk�0\�#�^�EC��FV��y��3~�{Q�:Ns��	|&�#,��$�^6��N9zo���-��i���S�� Cy8�E5�f��j^�)�@��a�k~�v�Ԝ3c��(�\t����3h3VF��
=�$�E��֋߃(cS8��42�O��M�ju��R��T�8˴|�"������q����o�Dn�IӍ�ڣ��+q�9$�<FN�_u�k�$�w8��]�@+I{y�D��u�L�/����Y��	
s�g�����I ��?{Z7����Hj�D���<K�'� ��ǜ؎
-�/%Gܘ)�gq҈d�L��{A	M�y`ԯ���_{$�rc�nG��)�F�T)��{���(c�I� �)kB�ޖ6���c�5�P�a�IS+�={����ؿ�'�W`=0�ôt�a����@��U�uԸТ8�[4��ʡj��ҋ���p=�l������f�=Z,�r[�Q���9C�{�V����)�CUG�Dd\T���@����S���l2d��m����v�[ ��C=ܶcz5�L-f��9�>8�;S�����܁����jt�����I9
�B"��;�Y5����p?�?��i�,����c)ʓ�S�,�x��S�Q����s�|%�7J��S�%�NI�eV-(�����}V��H���
*���Z#!ĺ VgH���V氲�\9��㢞���0�X���8��G|�����9,�)9�� u���oKPSA��7�G��'��XB����}냣�&�6��Ø}hQ��*���$9*��Cͺ�3h��#��������8�YU��w�?��hRQ9L��%��ƅM\'M�Cm�ϣ6���� `�4����_KU産G��,	���-�v���ω=���� c�����5�?h.��i���~�~XX[�_񓘳W�1ޚ�5=�Iy,N��p5���[#�0���\U�:;�J�p���g%�����%ȹo@~XB�%�u0���� ����"�}�����mBVE�r�BC�x#$U���*� �j�T��J`�q����im������[�'t"ͷ@�?��m;:��Z_�fK�-�ڿ�i�v'3��,O>u0��N�by?	��C��AЁ,�pg�����W5!�tm�k�3T�BYn�o\'ظp�����'� 33i��߆����Z ]��K�,5k�T�
�;�Fj���5�K�8!Wx��� '��RE5�ڨT��v�*<xb9xU��f��'`_[�9&=�!�� N�A��M�R�6�pA��?u��G�;5�S���j��U��I�`��s�&�/d4��$5%�XX�A��ϊr����;����r�ߴH@}ć5QO ���IzdU<݉�����Pm%{��q����ʥ%692zʈ�Ø$L����ӧk.q�mT�bm�'�f9���W���ޯ����l/���w��+	մt�G�t㡓Ps1������@�&�Fdm�%�D�A	�Bn�?�N&���5��?T0l��!Z�c�D�+���a�n�&�%tp�^��lৠH����T�Ud���>|i�:����u���F��b ��_�+ q�Z&��DD����Kp9^�����]IM^&�~V?h�Y���$��l�ϔh+_g�e���jYU�ۄ�\{+��	EI�W8�,�o�Wh����ჰ��$���5����OW7��H��Y� |B�=���'D˸kDث���9e-�\�7,��F�㨶��q�W��T�c�m�� <9���o�j���k<�y�I�F<��@�h�5#�zP	s;�����(���-�LR��3"��7�B�܍
�ek��0��D���7|ͺ4���o�9�.�FA�DQ�d�U�Қ�Y��8���q�z����>&G��z��f.ZRc���G,�.!����������dnr�������(.� ���"t=�|���aS��1����6�
K��B/��)#�+!fzi�5;;.O�t>��[c�X�����o�x5�2�$�Y+���^��dÅ���%�]�Nݻg&�^.��ٳ���ܑb%d�w�M��2y���';��j�nX���)zh��	'��5�'+���`pK��\{-qT��5�6׶��׻|A;zQ�a6���,��+����bJ�%^���$��n�5�R���)�R��&��'vC�c��x�U�1.���+m\dbE
F��\���\�3���U�?S�VRn���0P���|�K��^"�s��Y��d��Ǎ�nL�K�V������\�Q��B3��b�j(l"���hQ���e�C��a��C���Ltw*F3�fL��y̼��==K�P��J�o�[Q��:��O��������c�\D�Ψ������9"R7e�4vPd���3���f�1��Y�6��ѽ<���=rj`�KQ�p ʢ��������M-�, }���L��QVC�^��%՗�O��	'�C�9\8a�b�}4^�@i���+�ϩ��ߋ8�c5�)���2H���p�Ja:@��@H2�p��O9��h�Ù0�ߔ�2���p�N�r�j���\&�"�U�qk1��淟�_!�/d}T�N�z/�J��6rI/�##�m��y�Wv
�׾����h �p6�e�Y]�M"r��bw�v�;i-��I!dP�qe�����e��|��,�����X/@A>f~|v�j�8�u��~�����@N<bsI;��	��S��j���1=��L�W���ؐX��e��őX����c_�Xv-Wa��K��X�� �//j+�4z�US�W�LN��h�>�P'�t���(MYͩ��{F�bs_&^D��s��s��Qj�6V����{�d�Jk��g�)V`������M	��23��A���a����|�3�rR��<���Y�7bۺ4@����Iu��NTX~�H�'��]� %��'(�:����zr�ԯ�}��D&rߊ�y�
A��ng�['�l����2Fλ�pK�U-���)J����ƐzU�+س�/�f���&�F�Cp��+%2I<8�Ԫ�� �d�B����ZaV�I3�]l*�f��ṆS��>6������r�	@ݠ u"���K="�a���oA6��c���<��S��⠝��C���g���_��`�����%ā��30_�,!��Q��A�&鍴�ǔ�{�kH���m�߀�UWEεXv����2�U���O�"Z5DJ�7�o揼����W���vxl���Q���4�.�rYm܆@�����B���t�5d�K��9�Pf!��?�0*1=�}�i���i&��)Eg�v�o�
�0��Ϟ�
����}�������ɩZ�ϟ@H��B9�(.����Y�ؿoŸ���e]/BE�ML�3b��;������q�SV�Zy՘8���8'����:�w4K���{�;�Q���C���hg{����%h9�|5B��E�ޗ淵US)T���{�1���]ώ�&6��/%���|9��	)A���|)�%k����~A�=Pz04�JɢS�Ǉ�H����M�E�9�����G���g���D�K��<*�o*����nG�KR�w9�$~r��)�8�]�J��򔰥w%)���鿲jLYW��w�{2\�W��}�+7�+;��9��g�7	D�^�d�o	K%<H����j�5�E֤'�C�%=�������� �8� �����|��)��֛[�Ak^�9�����\'�R���~�L� ����uT.$��u�aX�7�h5Q|Z�m���`����Ł�r�Pmx9��s�y�q?(jK��z�#�vW�Y���4X�O���zPY(���F����j��#��H������/N�U0��U��*��({7��m�.�m��	'
J��%^r�0�o�s�C�[�y�^�V#�Jz蒬�2��������T�Q�_��W�I���I{Z���X��< �F����4nO�7	]��8	�֥�i]\9u�'
B�� ���F8W?D��8)�Д��l��L2�w�ǂLZyk,�̼�X��>�G[(����=��	o`�g�,�����R�H�%`�-�p�!R�Wn�0�*�קb�E�BY�c�wD�9���D���tГ�b�/6
�ϡ�ؔ����׊[#�Xp1K(J��*�k��[ 0�~ب��P��lV�F�4y���N[�A6����L��]���>]{~T�Mj!��^ǫ�m\�a���V|B�O��L>��~�"�o��m:*�q���pX�����w*���ϰ^����8�ι��ɬӁ3eq+����� @��#��?�'��,!�_��/�(�-�q����m�?��-I�J�-{Zn���hWŏF:�?J�8�o�\]�
�'��3�IY�<V_��#���vGD��@Ú�m��ETg�QX6���K�7�'_�*~�������Zփ���Vֲ�]�����Tb�_�>�|�!TZ�B6?X�<��vژ�I-S }L�]!�u���6������P���(y��l�TX���la�m�ͨ���I��q�qS�t.���Z�m�?�3Ѣ| �ǿLW�cJ=��c�=e\��KG�HU�#��Xu��W�ӌ�Vއ��CTP#x�m��FT��C/��]X�r���XE�{-f@2*�">8�5ol:�+�;H9Ն��;7O�Q�j8i�kb|8�(+�)�6��e���AqQ�?��^�pv��#��9o��ݱ�@���e�H˶��9(d�V
O�����!�J��8�b؍�I	��f���'�r;�;_\�+a���ɬ��S��F�Z�[~>�n*YZ��Ԩ���M+���Pu�\��@S��n-�Q����I?�sL����Q��=�Z�RJ���1`�Yv$2�X{���dQ�M�䅕�8��^원ȼ�,7uwҺ�> ��w0���9�+�̔�kd8ƿ�uOZ�lUؚ�b��J��kc�;�!ܖ�zO��9=Ռ��ѿt|��ۇvY����GV3��8�"')my�.���S2��h�R�Rm�zLպ����4𔺠 H�>,�*F��Fh��%�aΔ�D��_fUH�e#��N�w��֓q��;=�vQaask�
u^W���l
����%�:�ϻYq��K���Ie˂���)�����%<n���yF?��?C��d9�7�<^�I��+��$�V;L�-\)%x����nا�ˆ�?'9�a��sB[�4���6Ф¥[���ℬ�R'��5汔Y�t{�[B��#&���F��u�oT�P������B���-���_)���놫����~ 3�_ !JY�Ts�������kM�e{�|�"�W�[�}JL�}g�{�D�K�bߴE]��B�� ���	0�K!���Wv�FZ�d���.SBh���[�7;����i�����zҪq��C٢������.uO��xw�< c�rX��G\Z�� �&����w�י��j$�A��o�����(�om� VXЉ �J�~�- jlѮ���`�~�
�#��E�ڃؾ��}���Kݸe�w��:�>[������KP�48�ML-��多�1�F�0Y-z����1F�hY����yva�I�>2H�0h�tJ-�S�A�]�7(_;l��H��y�dX>{�o�C{���W��"�ٕ:�7�=n�F]��a�bʚ�wcdݐ��3�Ft��7p��q$�\���3a�j�a�g�]����,W�v�O���4�͟�:��[p�� �wG1�y�;���U���~V@�^�^>�k�Y�{h�z���v�TNY��
DP��a#��:[�^(VZ�%�O\�
�@S��A[�"2Km���ħ�������yEc��Ky��`�xK��� n��z!�3���������)���� ml��{w�����V����NF")DBn�e�~��/r��B�ӵ� 8w��4�(�g���� lfe��n��R�U�*�[)��m�{����OV��p�up$�:����h2؉�bL�y��nl��\3�������W߿T�/��}����j�l���Z�G��#,��͛5�S����d���!�P��uï�(���χܐO�	}�s�t�#@�Yt4�'�)�ѐ�G�Lo�@�#����ᓀ���>-E�1�Z��� �,���V1�`��O�EeW�g�"�d�w�u����+�l���G�]E���yv����6��Cc���M�@��<����<�Z@��%[�2nkb|��ǌ���귃㈅�K�_f9�W�]�����H�i���uߥk#��>l�u�6j��=�����o��%�}��|}��`���7>Ok����R����P-�%�ɽa�a��3\�P����}�-v͗�>���b�Є�g����|���6[��-�p���i�S�_Q�G��,׸'�6o���(��=f}�Zʹ!�t�p��-`�����a�Q?�	���rK� ޣ��O�[.jZ���3�$�K���#!�/8yB�MK�	�8�_�)��G&��g�u�	?�3j�I��i}��&�ro�Z����t���K�e�����tF},]�8A�nH(���Z,�E[�em�K� lO�n��ϟL\�T�_��2;9����A��V��E��P,�p\3��w���xF�Q�@%SD��!���&ҝ���5��F{��t�������عT��]��D{����{j�*��f�+0�܀3xG��S++'N��'�7�{� ��0B�Y:�mJ�,�wV��
�v̲1%"!�<WZϻ�|R������lO���'�-쏄t������ϳ(k��,�~@7{��1�|�����K��k�%(�:g~����ϓV�8`dhBfں�^�X�S��1���(�����PXX��z�Y[G������WJ+���YQ��j�����|��lCu�^�������G����*�#�_��R�Þ��t�����lo�1(�OP"��b]�������EG�a�Q�	w��xI��7����'v�V���p3�a|x0�/�� e	y�n�k�H��
vi��.��1@�z��-�蛴�燐Ζ��j�G�bs����7и����ϵ�ɧ��KzgG�����lc5�$���Yf��BB�d����b� ����A�� ��Wz��~!f�*�	:����rS�a� (��|H���@U"C~�'���d�Q�������[e�j�BA{���G�f�>Ƃ��P!<�a�9$x\R��)*��s��4��\�����/�8�&m�v�I��r���-�o����s��{��HÑ�¥�/�"���~��E�%�<+�{]��>e�|��{�D�q�z^� ���[{�1C|��#���b��B��d�h8�9��c6G����أ�|��R������/\Q��k�(�H�yE&ALo�m�ۜWP��F*�Aդ
a׻A-���Q7��]��T�qi�M
,Wf��	�A	(��r�C�����ɢk��/��;pN[�B�¾�C]S��x��[k	j��'NC}D��FjZ�o���9C�9�ڀtyN��Y��J��E����6�� uߒQ
NqRlLڸ�����OQy��(ߧd��?-��i���X��a :���`|��;	�݆�36q-����d�T��[N]���1-�G�o0��t���I�qY7/义�39�����u���|̮�r6��هܺ����:\Y9�axs: ���^g����� ��I�q�&Α�����+��Zd?��Sa�L`���A�l0t.����<��LH͠��e(�4H)�m?��7���ܲ��Ʈc+ ��^��ie���Ldx�Ukv�wV��8<����/K�_+	��*�<0��� ����`}EK<Ӹ���晅����XFD'���>��<Y�
Lb����Ǝ7P �l�/�5�md�"kz��C�ݸ1�4�n��ֶ�8ǂ�et�.��?st���,��91;͓�MĦl�~���zT��GC��$y���Ff4�s?G0;1�Pr.o��i�CF���YnXt�Wd}	��##6�1@]�JL�ðt@��F��! j�J��%CȪ��b� ����)b�&D_����ԁp����|:�����#�XJId�$o��2c�G����;�E�OWn���O��x��ݧp*����&�
{;�r�_�o�Sq�t����|?>ϑ��F�G��[ȓ;���5j����;��-.tՑ�;�t�S �ݮ{҈}|�{
q5�1�k��g�1(/�̦��*�B�`��Q�,�!���6ˢ�|��)[j.|2��z�q��1WZA�����7��_1�47z��, {R5
�[P]�l���K�{����H�{@�q�6��W��M�B'���r������s�ٹ�dѹ���8�!���o��Ϩs�~��y�/�	Mey,��n\'��]��{�x@[N�ST�{��O$.�JbX^v%���k~�߀� �FET\e��*��E{�T?�?/�9�n�=#.aQ���e�<�w�~D�S1�pa�����<���Yz��c����7M��՞��s��j� a��E}d	�H�<p!�eY�>���i7+�X*�B0�<p���l�-��C��/�ݏ6��a$SX���4�5�������,M��	a�[�B��ʫ\�dB~	�\t�(�Ś�,lt���}���;0~�P�)F/�iJ~G��8���S��"�xs��릔Ae�s���bz�Yܜk���*���Vx�40��<v]=
Q���0����Mym��i��HW/F��&�9w���F�=�/�2�Rk ONi1*�-����_��o�z�~���d���bΫ2�c�ڛ�Q�UZ�[>n<o�R�*<,'���OH�}!�<@|�^�;{?~ ���LЫ��w:M�8V ,����l�7��q�?b��='�ɴ�-b&���L�$��ԫ��6^�;�D��Dj��?"�
	���#���˙ �����!���|�s+C1�k"�@�t�u�a��-�x�T�%���,�l�{��H_<W�Vt��C�An���4�l�Ex�����_�t-��O5� `)c9Z�D�d��8K7����2�ji׿���t]�F��+���x���vv�1,�����$V��V_��-��n�e�N;�T�k"���o���j�㗟��eY; R)�u4�<�K��~_d�]���J�
Z�+uȎ2�����<�Ǫ��0�-7�ӣ�$A�ؔ
�?hxU3 �p\qd���=ڡ��,�c=���4?��~4}�ݪ#�;��8c��w�"7Ok���Q��6c[�ޘ1���K)y�%����W\� \w��p"@;0�q�E�E�ƾmTW�w[��~L��4ߟ��)�R�	J��S;�sV�zz��GM}1�q=G��K��w�KW�p׶��DP��[}�no�6�,���=/K�v*.Pjo��5	[�T=���MU�"^/�;���f�*`(Τ*W̚@���=�|4���*G>&&�`�WE�9�0� 6�~��7eYj����-N����3N�mZ_H�����`�tl������Z+)�����˲�lJP��/=maɯ����(�� ����8z� �J���+ ��ߴ7*�����aXp:.q��cf8���|"�fz�����OD�<���O�ɋ=#�:\� �#!���Bd�u,BR� �X^�������+֣$��e)*�8�lm�ޮg��["��ǹ�}����z����|떆C݊�¬�� ��ɗJ���[F�IM!* �9;�ON+8�@q�a?�(�E}����c��
ؑZ_�LYӈ(x�5� J�Q7�M���p��V�E�퉛;r3]K��l�`N�3(+��mW+���[,f
ʃ��մS�:��D�����%�M�P�_
d�'I�C�sb�
��SNl�/�"���5`�֕�����@�Y[�yܟZ����p� �uk�9M�Z�������M�l�
:��I�9�%&��"6l����ح] ��'�v��i7���~�F<PԿ�o��I:�@D�7�%	֋�w�^�<��,�D�N[Q��;'���W�I��?��_z����=��<��D��? w!���z�B�Y�z��|UJ�^/�)����~r���g����ֺ6`�J�3���hj�Y�������ϟ�]������*�5����&Ѫ0�]3�CGH��2cq(�����\XNL�\u7jێu�<�c���ŏ��V�����1���T'�$��5�du~p��R+�"��fDV$?���_s���^�;f��� �l�	{�겗�6U�m��䎚��݈[�&�i��������ض:*����ID8�|c𙍶� D]w��T����Ϳ �.������a�A9o�S�F��I����2���Zڶ ����Y���h=�HO�/��ZhP�����2s�8@�K�ӡ|��t)�(2��M�;�π���ܖ^��pz�j1۴���<�䜭[��_}0SE�S�������v��E�*j��T�kK�<ԝ��V����-�ΆA�``g٪4KHd�Idh�X��0�&�Z�#����K~��]���_�c�g\R���lRm��˦��4�r���*���P��K�U��r�,���ѾԴ�ˏ:X�#5�-�&	�2�a�lci�	N�	�3=,�"�o*���}ڞ��1�{�����_ ���T�����[^�t�1�5�-[�b�`x?P+$Y��6�Oֶ��.:@l�sfh��$8�����{C}�Zo8�˘�8����	'MJM2$^���љ �Ь��gv0�������q�B���\�`W��ѱ�*�>��xT��N��YGT���_A&�mC��-ZÒ��U�H�w�2�iSlY�a$���1�+�9���<_'��c�w�b`r�I���5��1U�dYh�a���OGH���c0$���7q��RBu��IK����k���o5נ.j%��,��l���ߥ,��h5dM����)��&O�f�����U#Y,�f��+���W��+oa�;b�!6���� <�c�wUOJ�Mdy�ݢ�r2�@z��a�O��J����!�ރ���f]x�+|�z��?�����k{(Q'^�ީ����Fe4d�i@��ʃ󅇆�"�(r�||C�./O������?�4}qW	wh^�S��_���䠕y���s���@�)#�x
hb�Y!�f�������0;w�4�Y�A.<~���_&Gd���ʱ��v]q���K;��z���>�dZ��eWD��+�q@���O(��e�F.ԭpf���K��`�dYU!?���0 U��	:-f��
6ja�oM<��71�?,Μ��C(Ҿ�Uw��QFux�8.�[���ԑ����<+�L��;IIřN�ݧ�2w}&KQ�܊%c�a������$��{�B[$5��쀗��\��|uTe4�vmz���1 ��$8�n�2�$_���|��2�e���ހ��a��l٭����ٿ͒O@��)T�U@���zȹ�9����h�[�����mt-6 �w�{~ٕd-:��{���}��;�56~ ���n�rC�dh���>�������Q&̩�[|1�"���r��,U��f���,��/{�w$b��g!��L6�]�^�:͟�_QdEV/ 8T�D�Uj�����ʲ��x?V4�f&)B�R±�Th��P�t��D�G�� }��e���Hc ��]�aW��Et�`&�Bq��� hi���-V �j�@O��0��7���UrLXG���0���ۀ��:����e�}Ij�i�3��1�D�������a�lӦ�Sxt7��ݙ��J
pUw�AW駈>�E���k�q���oKٽQ�o�ǰ,���$�� �b5��,�P�'N4I�j�I�m�x�`x�/�̀?8W�}�Qf<�.Ƃz����[�k��_��xuN�2{�kr��n�r�V����+М����'p~�-��yj��|Lia�K��l��wpqHw�<����YEBq/K�y���&�Xߊ/O��`��!�^�Bd��ڝjl���w�kms��f�	E:?����ip�8���Tz@b'�1������������*=j\���p��T89���ſ!�(5�_������[Ɇ����j��_��7F��%	�ց���βC<$�m��q�D,G�(9�0��,��~���z�
�JJnlƏx�Zw�a�桬��wN(o�
W�ʦ�>&	+歉�O�b�@9�����O�j���VG4�E�E�v��sY��4Z~)t�]�>g{�uYP��Iu�-g�q���������<1
����#~F�\��O�2k~�%Q��oé�t� ����w�<f�����lߑ�aSH]�?�?��?�YH����9nٝ3�-�����k����Yj4�Z�[���Amp�P��^&&F,�9"e�� ������s��"%N�ܙ�N7��k��(M	}��&Q9�\A�ض�֘���|rG�y�o�_Ѱ�[�m�C���_�u,��WT�)��e��*pol|b����۩>���p�T���c������J�&��^ثƑr�� �-R	�߿��+;יT%�l_w>���R�*��	V�#�%S�&َ�0��ҧc%Y�t��W������~�����J[7�Dn%u�sX ��$Ӭ��mU�c�_i齭c^��kn ����w`�<r��	|��Y��q��S�Zs�!/{M�./6I2�����D����Zk\��}F���3L|���4�&_����FBf*�۹����ҭa�4��<��A5��Y	~�Y6 ��Jޱ���YA�(�b����)��� ��D�m�໾O&������hmf�ŀ0 �	^lR^�-W�;K������9�Z��r�l�e[E�p��n#�D%	Ǯ��¤ۜ5Ͳb�;��9�̙��3�B����g�����@檧�7�n?^�v�p���<6}㇆�j��C�E�%LN��)�u��sM�H��	�s-�6�H���
Ab.&o����w�ڟ�Z�s�6V��kֿ��]
�o�:}]U{����NR��jK�9�PB��4�6>��W���mG�)7��5-��z`@h��ľ^eS����W�39ҍ���N��&;��|� NL��J{Ŝ�@���aE��e,?����Y8"�\��W>����Y�&j�q�wpk��ÌkMx!i�
"�b���Eh�Y}m����o���>U��$��׌�?�^���2�[�a+\X�+@�if�붌H�b�@� ��#����䐜%�R�L���;���M��ԭ/�D*���y��(��;�>��Ta�^�)^qA�.;ߗQIH� WG���ÒIʐ�8E0+"`3r	�*���:f��,��UЭ0��,0# ��*��';�G��9 �;8�D�@5ҭu��طV=�}�XE��V(�$9v55v�m�c��g$�f��X���z�FmOU1c����]�<<&���Gs_����2��Es��K)�@��dn�=Z�&��tj��x
:js8�9�(z!�Sc����eC�r��{�&�Zh.�Ð$�r��lTL��?ɘn��cB��:�F�t@�]Mh*��HOaG��:g7�j�����BЂ����AY���!��� ?����_������} rd ����(�%�{�]�Z��ݲ�VN�ҲW@$���OTL�V O{�,���lI��j��r��g���2��f��[��v��ć$��d�q><{�c\wY@�"�@),��V�Ҕ%�;�1�&'?(���o�H��А�ȊW�H��.A5�UI��9���3�ǃ�,�����^��r�¥XZ\O��	f��&s����i�X��V@tl�"�c�e\oq^܌�}qkk��=�[P
�3��t��@��Qx�b&V�No��s�O�x9U�Tp`���������$����G�m�[��*i�l�W�s(�GYV\>mA Oũԛ��.Ï��W6�\�t|H����@ݦ��F�TJ���3x�_�z�q���FZ]�W���#��H��Y��Y��VIR�����Fj��*�tW�~���~ly��з����U'*��YZb'J`b��-	���������%;�������g�i���}�������1x��P�d冎e$eN�1���C��!��ן'�Ѷ�'��u�@o4��lbC����Hp���4���ֆ�(Yr2�Z[sm���B�P/VNez����M=�o,��$�r������D�"�?��
��3���"����l|	U܉�@����3�������$�$��9^=4�	��B~��.���|^��UX� ��?����1�J b@W\)1�qa$u��r�`Ǖt�"R��6<&}��Ψ+:��7��R�����k���	?V�Ћ���P�VɎ�m���+��8S�i��V�x[wyx��9A������Bc��iY��M#6-�8
B��L�~�Wse:L�;rP|�2��I�G�QB�T����A�Z.W�����_w�l{��Ո�Z�V�,Kfl̫C�B�RW���+��"}P_�G������y,�>���x&��'�x=��
�Ї�W'��t���,ѷԼЙuUT�\eԮ�������~䫽���y/��Fw�uS���X��i���J��1&�����8�FZ��F��I��ò���Mn������_��G-T����$8 �IUL�G���|���H�\O7�>�j%��DB�U���b4��0��Cc�K��Z<S�R�Mo��{����-�2$S@�v}mr�tXK����i)=K����A��Aܙw� >�.�Q������Z%(5��4hFb�S���32J��٤�Pc���zڹ,Rf�xsg��q5��=%�32�A���_�s~�A3����U}���y!�w�G��GX����H�R㍉\v�k��o,�#~��0[��F+z��k��;g�������4l�3��5f��@�f��:eIخ;������{��"�
I�7���P�N2b*��x��D0��m�=�8���"�/6�|��1�Z����ʫ
���O/H�s6�#�=u|�;�s�	Gf�������������Һ �.�/�*�]6Unw.�Lڇ���!!�voxY�n;�#��(j���2�Z�s�Y���t�Dh.����T(��C��ճ��X�?���#��v�NAD#Fd������W��)���
8�J}寎�>��ر��(��8�^B�R6)j�<C�N^8fQ���AX.gº�<�����I�I�lm��I�Q�]�'���FY���9b3ҽ�B%��]���aՇ��]�Z�Q($�^���������ڒ��Ŧ h@�&�~ �j����:��Nf��E�ȕY���!���Y�2���ac�k6&��v��o��N��6��!;J��3o���[���k"���d�X̂��[��:�퇟A��1mQ3a�7�'F�\8T�`�0���\�c���k��ث=��1����}8�ڳU��\Γ�g$9����}�E������B��ՔK�v��B0����U�F�����x�Z���I5���a�Խk_�
a�s�gkN̉�܌.�Mk��S7�@��%��d#���MU�[ʆ�Ny�Q��ߠ�)�N0��$s����"[P���r!�����o=s~GHM�T���g��q���ӝqrƍX��`��^:�%S�����t�S.��,�+����
������݃+��s�97��vkD�p�v����$3�!Lt��\}����1~���E`p�m[B�trm,�n|#���)��K_?�Y����y�l��R׾a]����Ŝ���V����;)n�9� ���y#B��ǰTd�8�{H���yc1���o�5&�Jn^^��&����&�%}��6�y�`��Uz]0\q.#x��y�'�fC�\҇�,ޕl����"p�F��#�Cm<����"����D�8ov"zț܌�08M(�&j���r��p	��)����<BN��[���*��=l����daTO�N�����ʑ��������>���qT�?Q�(������� mKE�8xZ�zW�7�ɭ��&��s�|���+���zS�B$m�A���r@�\�s$0n��}����oRZ�4:�L�[�=��~�u���]�]C4�w"u�}tHM���NS|. 07P|gAX�B��M�>���^h�H��{���(	�Sq{�4����o�uvmS��G�my�A@���pf��ɠ���ψX����6���+� �<�VK�C;��x7�z�<��&x�Bp�ܳ\\�~c���W���)wP��aK=��>�!|W�����Nـ���=�(^B����}⛸4�w��֫�˒���3EkӓT���I���hЅsiEv̎�LG$'�e'I�5v��*/�	w�������*�R�`�n��Wq9�TN�fzhFȇ~�7�������5�Q����J�e��2��č����;5t��vZ�R�_�u�ƫ���4����5o�ӏ�f'�T���1
%{�́hח,�8��^�wˤb�#!��,⃱�"�����)-����S��U1���F�@C�tgj��v!$�b!.�o����gQ�I���̋��3�g�?J�-b�K���BWz�1W�ֲ0�n.���Vb����LO�W�m3���;*�ۆ��m���B�L�H�b�Q�R�7�����,ovg:��n\{�(u�@�9���Y���T� ���*�ٴ���K�m�� �H�CotVC!���G�Z�j֌Q�DBW�zl�O�$���P���7^H�n���2`U+T��7�/c�c-_����T�.KK����_�����g3V�O(YYk:h�<�M�f�! ˂����hr�0bX��I�J�����GH�ޟO"0yڲ�T��e�t�A<�3퀵�:>*j�*�N:,S�m�s��Y �-ɽ�Pb�갇������<Yx�q�˂GK�_Na-P�,��X/D�Z]�L^.1g���L��C�9/a��@s��O��l��=�6��?0��+术$�YA'FpZH���E\\	!�PV<_�p����(q'�VA��"���;����{������h|8�*׹d�~�����R���p�k������BR�^����՘na�q���v����@2!�7�p���˺q�_�8�$�?�J\��=��?;���۴"��{]P�LW�1da����f�_�&�BK���k�I����kd�~h����5��f5����]���O��v���ʓ-{m�S���v>��V{��)�0����u�V��8�e�� �I������<��<��r�m�C喳Á����y�LD1�$k����J�o�P"~98�s�筦�� �"t�y�Td$�ޟ݆����W�nE� ,�
2�U%���?"����u<f�[i��M�*dACT�RU̯�8���-����>%�M�3E�"j*�65��_��Ͼ�?�e�i����x �_�(A���1�x�ÂX�IVn���d�m�%	8�	��/]ߐoV*q;��U���n����$��k����-J��#Ũ]t]����u��:����OC���AQ�O�}3(Y��J��lF���#҆A��x2ؑ\�Kd|���4U_n�9����FgOR!�p�0��j��FB�0ϵ�k���Dj����JVR�P	%� M�p�p�s�����v��Q�̡o{���VɽO^Y���&x`9�����������A�0����NK�p�OXɘ�e[y�D��Q�8�c#O��6��9�F�t'�N�'yՏJ\l��yK7FW��"��"dg�.R����Q����9��l'S�#E��r��ғEBz��{a�9��~h�e�y�?�J�C��ў��hyB'WK���9�����e����
����s`���_�XZO�5F���a|��2�3C`�/����C�x�R�MCΘg�aͧ�e��y��{C��=ڇ��it^��5dG�H�He�9�Z�w+��k��F�k�|Ǒj��w�b.�ck	�z��Z���غ��ln@�=G{r@P^�h8���5�[��U�
�H�;;��Э4V���]��"xZw"]�	KX��;͞D�����4�����>����z�K������s�;~���]T/����i�v6i8�\c��)m?��p8l��
~%���?&�(��6y=�Dqm��mY(Y6��R�����q@��o�<ǻb��)2��c��6T�ʌ��jb��CF#���{����U�Tm��|��,����$�`W^I(��Y�:ԛ�F�˞�_<E����eH*�O��rg�J��b�rAř���r��>k>��~Ȧ���O-K�dO4�y9	�oT���R�)��F�|F������K�����{�],���	m��+(:*����0�y5>g nA�Z���l�9y<�,�źT�s���ܔ@A�+B�^'�8I
����f]�kf3;4{e�rq<�����Q&�U���Gd[y��g�Br��@�I,#@/�Ic�� �6+<m�uZ��g�"��5�:�
�ϕh��Ү�s	>W ��HOI^-{W8״��M�D�<�O�섐��\SC��.��m@�6�1�!ơ{u�\I�����u�//�TU���gV��tgz�(�#|,��S�^����P{@�񁄾��,�1�3\�O�ϐ�b�g)����Ӡs�嵀c��)П������s����X��J��i�Eˎ�bt@��JV�LJ���sXC���0���U�O�1�;@Pl�>�(�ʖ�\�0���0�ԟ�<t\�In/���*8k�U������1���u��{���/��Ukw�Z�hǆ4aG��	��!�a�N���L�_�d��D���v�ΟOo]z�Z���Y���o7D�`'��>E�.q�;�Eް_��hB��^�0^5������х�!(�'�2l����^��xW:�8R�<��P�K7,'�>4Ǳ���-s���ckV���-�H�&N��d<���� �ʌ����B�`K�Ў ���/Uܖ���Ӓ`��E[�n��ru���<��/w�"c���4>��x���S|��"pܞ��݄���I���_�r�!2_��A�H����(����c��j�'��m��B�}��w���ghHA'^���--Zy�x�������Rw,��I�W�uo��6\R=���^��.wV��@0��%\�q!����|8-���0��p�C � a�8�P��`��h�\�x���jCu����`��h��)�%O6�|�	Wl��2�Q��
��f�\(D�,����LL*2G�s�P���C�ʀ�rEk�Uн����<�`�b�چv�1�Q�a��#P^����XA2�3T?�/���L����VH�(�St��=i7��O��Qb�l�ϡ:L�-���u٫�T���Ni�OZ�ևk���實8D�ٽцT���%�~�L�xx�����sppXR�R��Ǫvt�JSNx!�6\�1ʘ�O��L�����/A�>~�M{ Gb=@N��ТǲM?n7ۭ��2��6�m~�����ҋ_�t�g:��$��[��t�	�\\4�d��L(�˸6�
_Q?��Z�Z�'y0�����>ןTG�������s��0G���w�v�?�G�o>���ʉ���-�!�Y�체c/��ٮNV$Z����(I3�
��f�x�V@N��^��X���,�{D�N�v���]Ķ_��1�;�[{B� I;j�X�)jP���0��(�����rz�^�jf��о�q(��((ߎt��>�7I��-���k�qq^q- ����$}�����[�g �1�f�q8�>t�7�V录���5�Ք�5��:�c�/��sM���F1�u����6;٘��$"9��y���0p���[%��'�~���&��I�c�tPy�d?�H��>��9�:�[}s�bK?������\��]�v�6��'����H�p�LQ�iM_'���vL*.�˔.%<��;�L���2ςk�Ÿg�}u<M[���E�{?CSe�*�{�qXA���
$��=б�;Su�o/ájV�16�R�N��	�7�U�ݠ�"jr}���nw�iB����?��_�Yߨ�?���xJ��c�	���Ec�� ��e���,@����|H�R��$���Ϝ��Ȥ]�0��̃h�L�3 /9ip&;�0���O���Rz��!(s�:�ژ"&�!{P�xE;Ծ���m��j�Bπ���2���7��*��^hS����Q]���w�$�l�����F�qJ�����/�F-B�Q!����(ٱֹ�Ϛ��|���_[��&��|�JX�����`�X1m�z��w�mN�5�<vs���Ixf��7�y1�w\�)~�`Ҝ׵��P��� ~�橕�g��� H1���I�r�\>�ԫ�57* 	�G��>��`>�
ϣ�֏O�&|���U+�Y?ro]�}rj5f��N}�%��*��y�8��v 
����C(s�b�#�A�:��Hō�F�ٙ���ɴG���I'�����8y@�����1T�(x�d��=�b��{�'^�N�c�!�73vM�%(@I��^@�"A� h�V�ngl�[� �k��e���8���0����r�0`��f.ϐ-�Q:0���ٹ��Ab/1����嘘�C6��7Ȩ�/�3r��bo�<�1��?��T�ӔL<�(�ٸ�]�Na�ԟB&;���:�E��o�b��*/sW�{�*hR=V����_�e#�f*J��&�(p����'}�a����٭��ջ�AEД���)����պ|�ϛp).�C4%q��>���[�!�*w����i.+ D��?�S��{��!�O�G�~,n�U�>�Y�
l2���vW晃��*	6�O�^3%� j��s��8��e�]��u�y4�\	O���́��V�>~3�d�Y�($���9@�k={��b��7� �lEW��s�v0����$L�a���~�8�-Jm&�Q�Mذ��'c�)����%��=&Jh�K��0��]�j�d�~�b=AsҎ��\iEθgJ/����&5�
�to���v��<���';�`�d�s��	���72Ĳ�S��\S���_��D#G;�U�d�C�"�W��D�*���7� ݸ ��+n9ca�dT����-�0���d2)�����(��*���ۿ�n��Q���(x&�M<�mk���߇[�A�F̈́�.��/�0�	Ǒ�(A¼�`��׍�;!�0,��/)ӽ��\O��{L{
`x�\!�`M����2�����eפ=�Y{�o�{YW,������0���w��Z��v1RD�H�0DTQ�
���q�*���:�����qcR�ح�1�.��,M���a�wC����}c[f,��/C�t
K�)�[r�b�����N�_=o�E��`=������=Z�r�">�R7xЋ@��پ��u
AV��)z�H�z�1�wJ�FNL�=�����8�~ ���(�q�ּ�4���E�)� ��Gi��D���3%5�f?�8)��T�!綡�ON�Ǣ��͙�,�D�(��;��
�wt���$�_�`�[�UZ�Ҧ��fK@a��v�w(o��'ގq��K�,�~oD�&baO��ے��:w��:�扁S��T�8ױ�����{�č-�?�����r�;��20 O�-�^i�3.�ɖul#��k���*vڔ��R� ٞ�C&�o�DZPV�1�7R��g��䢸41Y���X+K��i���́
����)�e�nv�EK���d&P���d�6�f�x��-w���li��[D����	� P�����?y5b��0�o�v��b�0 ��^O�E�3p�����p���Zp!�c<#C:D������vD8����!V��xS �hR�B�	&(��kz���6��TMq����d.�RT�$��>��� 媼b�a�f�.k�x��%��lmWˡ���eQ��%Լ-YФ�g�InGm�D	��*M(.�?�$bI	z(��>op��v�dF^�(%��B�9�M���X�,<��u��ʇ�qO�G�֝}B�gC��H���;5ٍ��ɡM�;���<M�Z�9:<�yi(v�w{�c$���R��Q�R]hμe�Q&��۝�5�5�eF5�
�oC��y��~�1˲��S�����{�)�g_������`ldf���!J0p�<�d���O����\�w 4{{�����{��6��zF�c�a���� ]��*
 �I>uܜ��S�
���Nu�t W/0��_N����b���r"�e���*C��I�7�S��r���������d����������s8=�����د0�__���JX�q;���a*:��zG��JK�e�dۇ	)�s�}BiĬ�{b�������k���e�i�n��a�؄��T����e��)u�'(
��d�.�g��k����K�u�ڕ�o5�u fCі�yޖ�_\��o(��<�qZ�JC{�����oȀ��:��W����7�������lI*������ ��B/�l�g3��p�A��A��'�OB���\v����� ��������1�͑���<�c����	υ_�{t�lP(,�&���C	P)�T�'�&`b@�	�ISTG��v6��7������9����vVqЯ�4
b�W1P��0��L;u�( K��k������_�D��tH窬'^�:��w�t�K[Ӵ����#��&�ٓ>K��ʚ���ʎD3�I\:�������T[U�6PބY�_˖�$�P<Wu��E�>}m�@�n���mi�ctB́L@?7���ѾC	�+�ݰ���{�h�����)�w��7����h�M�ڱ�:	K��ej� EE��U�]��~J��/�cy���,hu�rDP��}�;!�_�n8�h�|Og�F�Ûzx)P�ʕ��u�+'`u�J��Ї�sDmegVp�#Ndo)�:s�q�()f@��h��m�'�ڤ��1����"�J.4�%��ь��+\�*X�W^�L�>8#�pok.ƊxVIhX�4#̉�bAx��_j���PE��<�8��� x�"�Z\)
%ZZ��2Ti�O�$r]BJ��k�NܖF���[z���PF8ӯ-��X���bľ���9~�!�J���i�3����ֵ������i�o�TX*|,�Fo���Pb��#�g��f�Jq���G�$�N�h)S�\�����X~�S2����c92n�G*ޗ��@�������Qk�D����(���� ����'�7�튠.��Gxpn��+���a�a\�K+u�4���R���J��~�T^WA$~�x�Y�H`M�F0�`*�%AF�3�\P���_���r]"?yBHi���;��2�2tt�>Z��� ��Ǔ^>�\���}��	�R	e�������Jt��#4����w>O��עh�!�Kl��j �L�<�~�c��G*�N#��a@Ìv�G����o J�Y[�`���@4�C��8�}�P,W������Ѿ�[=��J-����ՀՑ�E�2��`��n�"�P\(P@<��;Y��BqG�{�~H[M#�@j(�����ml��F	B�C�A��l��-�tq�zЖu��J����K���R����%��n?�|)o��7�}��(�~�r�TD#��Z�4\7�Z��GKξr�6��-�'�p�
=�S�f��o�yI�2�/^��ϼ��u�SlyH���!�n� x����ڇ�*�xz|�/�<f�Q�K����_ݺѲg.z�XA���.I���ʼ���W����ތ8�������Y�9�rhja��k�pc���
Gfn$tÉ�\���p�*�2sEX+$U����c�L�JՌCB٧]��|�D��5T�  �!��w�&���Ң���ا�4����v�jv��Ťoyu�X��[�o&gB�E�^�����N-�1%���I����n? ���GJ%;���Sw\]`���0^{6��ugN��H��:c/�{Q��J���l�mHW+@�;{�@
�fv��b���M��S��ZJ<�0��LS̟x`b �)���q#��\$e�L'�]��Š8�Vt3R
�(�h�����|ZE���������33�)t؊��-#�,�����vO��'��0���.�~a&��gu�>O��l�=�ϡ���E�1�Z,$�e�\� e�o��A��N��DO/_k�%c�իD��q�Y5�vqL�Q���Me_��P⒁���>y�V�>�а��b'lf�\����?n]����լ��&�)P�e�����:�d�?S����ʒ����H͋�}�]��}����5�-��E'%y����8�,�`]��S����7ų$������[E��4���j{�"��ʑ\��8�	���{lfp��`���0�B>Gn&��-��+�@����%�C���%��i͡�1�:�>eN�(����7lJYtm�%�C��b։g��E���Q�j���nQ�	��t	Yt#�e����!��	�q�C[����P͜D�]aק]�F�1�f!��l�t�,�P�<k������4��M$$�y���O�"J:lW[uN"Χl+�A�u�ʭ��Z�����g8�B�������}�&zB���h��X�Q�wV�a�B��#vMep=�.�K��������^��*�.���������k��U(x?hE�ʴ��k�"�(��C������,ĎLrk�����0w
-vA�捰�>��,6a�P}���%@���U���w�-����/�#2�3�����&]<Ď�eǿ��2s�,��`y���mb���^J�� ��6^k�)�4�ud@*��c+�W�W4g����ۥ�A=@�=�j�;�d&{�:Ȍƒ;��B;��k��&��-�����9���X;_�N"\0��	�#����:,�m V������>"�<,���j�W����2�nð�m�����㻣d*��8׳�c�G�)���X�z��$XDoV-�ZӬx���R(����☔��UqEK�ͤP��k�X��/X���'����hi��\�o�B�Z�k�HL�m��
�>�Q�(���ᜪv�/���o�Kޒ�Б�0�ܻ6�+�o��/by-�rUE�k~.�R?#Kћӛ�8E�`��Q�&�y4t��XU��ףrQ�����H�(��k4���Ba^̵�(aS�o�Ѫ�`�k7(�h,٦Jϊ�v�[�n����ɚb;�E:Ы{bf��Yc٪-N�	���,����M>�'�����Q��ܕ1�s���J:rn;�$l��U}܅Y�`x��
]�Bkk~�"�a����_	N�p=|�IuEw�{�h�`�%x2;��|l�P����r�$�����]8��=��]5u�쁽��~/t ٻ�D=�U5�=�B0�˿�ͼ��c�a7e�e�
'-v�����$�8��ŧ"������,rKy"�\{
���qCʧ�y:g���������� y+�`��IZS����!�8q3�eJ�*�
	R
1 �/��:�@�
rs�	!�$��?��87�T��D�C��̚sژ�0��d!-c/a0	@/� �����z�Z~�g�|�G\�f�hWI��nx'�c�K�ϴ'��6��N�����\2�Iz��-+*M�j˖���s��|6�|�j�W7�g�a� � ��ϒ6_?�Bh��m�+�ok�
�]��v�C[(�k��{wt�P��ܢ�H������|$���.�2H~_�l�o!�9~��n��'O��hT���E�O��W���`Y�q�*8��$|��EG�V�?SS�@L����$~#��P 4��z�o)��W���0:����
:���i{�!5X��26�w7Ul� $�~=v�u�65_
a��1G�����oC��=���zdzqn4�Ib�Q?�l��X5����7��� �f�vk��RU�\=�)��ӷ��5���$����HB~��R-���>O 0�V�!�༉p܈_|��(�%�jb�F�\�s��:�~��d�1M��ZB�<ٝ�h0�� ��q��~奫��-f���U�Xؖ�A��+�ºO��AKZ��VJa��9�\f������7��vd?�b0�;E�);��o[6"P�2뷅gk�E`�f*���j?��4�ny���9�����ߡS�J�z�Z�?�[a�i���@a���	8�ym:,-L�3�,@����B�J����s���|hK��"SUݞ���;a�Śث��p���j�U�J��r�m��)=抠c=$�=�+O�jM=�ĞH�����;g�F���81��	�$�Y��5\(UGx�O�ʿv}Y�&g�9�Y܅zX�,v�@�\���vu~ JdY����}*����m�-u;���ԙ6?gK�઩�����(�$����(哰	]h��&Id%<%���# ft�	V�(���͜��:f��(ƺ/��)�r�,ok�9b���GN1�Fg���\ݝ���ڦ29��
��H������:��L� )7/�݇�΁�P�l�K-�H7P���L��x�ka����U��D+Y~X�#�k�b��!Qڡz��,d>OǗ�h?��m�!IƚY��5�A ��=ҟ��L��-�\�=����r�˥-�v[h�HDfߖV�}�;M��QwL-[�qڂ�L�:���a�*/�����M��/�%	�i$	̷��WKKDȩ,I�I>�tĒ�1ｋgP�r~�C3iR1�S�M�8,�{�%s��s��Z������Nj�'8�=5�P�<�JZd��]9m��q����t�����O�Ɉ�
�U����e� _�}�(��S0��r��SKx�ӿ�����
��y:��Z��cU��,9'��)�F�(��š�I��<~���V���^h���<m�#�qK�Դ�w�J}��aW�55kx�-zJ.�i�4z�)�4�y=�c����7Y����r�YrIѓ|�m� ����{p3����J���O���R����t�R�1�X���>��������]
�D!�.JuȌ��x6tXu!7�i��f����S�]��q��Fҳ������,�uW p%Ȣ4�E���B���\p�^0V�7Wy;�®���_�d��:�ћ�u|!}�alҜ4�D;G��a�Zl��r#
���c�����Si�L9���j��O�������y����>j��V!��9@5����������q�ߕWE�g��JV��a���7�0����n2���YnL�����b�SjG�՜��l��(�w%6%�̙��S[:~�����I|��t#f�y+��
 �M���Aգ�-f�1n�5*���ʹ�%�Qڷ�A�y#3E̞�x/1�ds����X���%�J�V�*NR�7�Z�Ou��<8�gt�i�-%8#�P�'�	����!܅�/���V�>ț3N��sz��#�_Ԕ���> �;���k�����rw0�	��{|G@^��Ͷ�p��S�}�s����~l�X�7/1y��~�F�7w������>���/4�i��U���D���1{�����&�?�\+����BJ�iBy�<	yv���c^:���f!?w|;O||�p�F�+�%h�7T��@���xD?B+�-�!���lV"zj�-�i9�����J�e�5aUG��E�W��:>bPZ�������6;��$���P���`f�)M��vŦ2�W;���x�":CN,i�"1X�=p�]q"�H�*d1��0e���e��8�o){=U�͂#��j�fx$On�¯/X� 9!�pփ[��v
ʃ/�y��:7D�`�;�0U ����#�� HiY�N��U�"���H�&
T�#�<sti|k[�uZ(������o��P.��4+Sc�֎L���nz,��P���U�]4#2EJ�M�`	��P*(qG�$�(,'��8�%yH�����I����LM@r�K8��ܦ��2 w������u��]���@���P�&�$�o��m�ok!���YN��c�$[I�yXK@��^<���@������a$�{6�F�^�-��iO���q}���NX3�wo���7��X;��PKlV�{�Ҥ6�L��˧��GxS��W|����oб��i<�]��.S�[m���ccAb$�z�X���TP�I���s>�+���̃�I����9@�ow}��C� ��R	M*�',�v?M�w��=������ytF�OТ��3�U%:9�SUq���&1��W!�6ď�^��1A��<��6������U�E� �Ϲa%�6�|�@�L�[@���~�E�pVN��F͗���I�+�RU�f���,`�P���4d'О��%yy��ʃ@-o;�,�gj2A���&��B��B�̞�Y6����ں��� Fb�q�ޝ vi��{n����ёD���S/�a�F^)������P��{��ȳ���x����]�[
<��%p��2����gQ�q�b��z�a�5D��)��.U�h*8�n�w����s̻�a��x7-��+[�r!}#�Tw���X���M&߸��4&�_�0���pm�F
 d�<��ͬj�\�j�r����$�"�]�c�@��#�B�����E��aG�~�kL����V��|�I�v�
5�>��T;����P�p��V��0�(����,l�݂����%�)����nx�� ���Z�>����
�%m�CG��8���R�b�3�2B%Ђ�������.r�V!�G�����k��z�L��l���F�$dʲT�l
�� 	)�|�=4�!.�����Շ���}�?QE��v*!ܦb)�_�js̛��?˪V�$DB��!9e�W��5&��+z�4�BC���������=���,H\?k���OA�G��Ea�@hU~�U��QWy 4��zYy�(��������Sl�l���V\$��{/�d7��|_��c�O�<�l�z:a�gN��7�F�$��\\��b=�>������s��J��æ�&O�O踍sL�	��*�b�0=4�	O����	��au$�e/�g�[������Į��j5)omH�i0�ɻqQl4D��^?ṅ���>1��.W��R�d�FT��ɇ���W�)��kv��t�S�Y��gk�L'���
wU6��2�p�g���&��ϭ��N���0.߉�cf�_앣j��Dj3��k�e)i.k�@�I��/'����;�i�*��Rp"|�uӨ]���-Ų �?M2P��Rթ(�4/�������'����vd��x���0�y��񢴤�ؾ�3!��|�r�;N�U�*2�CO��o$B�/&4$�f�d�\y�V��_k��� ^Ypݧ��DآS�2,��]ٌћ������g�sb����$I|�{i���	s!�I��[~q��AUS��et]�>���2F��\1�2]�2SK��#�X!��>vω�e����Fb9_���p@3|���/;�܊&5^�mvRp�K�ꖃ���Z���E5\+ƹ���� �d�������e�������)�,�9���rkISQ�:�*J�����f�}�2@6����l�
�17��s���րM\�'��Q��&&�����{&�X��oѺ���v�iURE �;����Q��B;�l�<�_gj��$�����7{��v](���"Rt��h�3����n
&�eo�M]���F��\rHU�P �&a����CԮ���)�0��9�´�1�Oa����ޓ0<��|t#x�p���qC�{N�5a�28�@�~v1���^��5d�w�n^�nF]���%Y���e��e�z,�r��J�b-����ˁ���|-�y�6
p��������÷��%�L�Z���ݍ�1��e���ϩ����?XI�-�sX�q	Gj��&\����k� ��kN��_�\x���@�(FW��??���A�hڣ%g�qޢIF��*
���xߧq�Is5D��
������K��' ����<��t�ٝ�vLI�G��t�9��$򬗿�bt?*�O� ǫwd{_��.T403����e�LX;i����i���s2�?`�B�8�#w�*[�L���� �
�
�a<�w+6sU��ibZ�s:W����߯$2[0�	��Kd9�tϵ��Bq�4��f`��.VZ4eٽ��3������`9����	��w��޴!��i�\�(��6V�&�l����
�9"v"m�yBB��X�t�D�I���K�>9(�%Z����N���D1'�SIb�I)!<#��E�E��hp�1)V���%�i�'�*(�r���V�j���9^+�@ԫ��a_�b�5]i�Z�Ж"�����mИ������f.��*�B�)#�� �my���/�:����ဆ��eH{Z�?j�����c�ˀ$Q�g�����f�&G��^7�C���-�>ќn����ƭn��gd"�W5Q>*��ŕk�ӡi_�?���.�lg1��ɞ�	|�!�v�f�YU�/�$W�˄�i���BN��iߴ_V�	��Eܶ�Ds�U3���=]<�� u���Hਵ/*c��Zy:�c�u��'�D=p��7 �0��o����TF,�Ͷ��%��������!S~�^$4��U�B�q,=��</e�61����"�$y?���h%L�a�hg�����5#���	�Sl��i`'Wҝ?c��M�m;@�;����},v�7���ɴ$,����X����	0�����c�ǫ�~����5T�qq���<��ĩO��5��8C�������S~���3���?
�j�7M�`]6f��+[�}��5���9��.�v@w	߭5�AH'�n��-Y>��{��Z�~�<��5����E�:%�n3��/�z�1na|pw����8��u�K怹��z?d-�UT#��s�6Ĥ���3k<-AR��7f3Zj+#���4��˷�&O|��
*̵��O��p0b����i+.�m_�����`g��N�:��K�ie����g�%�'��y�Lh�V���m�n��a#�D���ԕ|Ig�$�qӄU�RRu����gK��s���3��u�����y�{Kg��g�}"Gq��G{pU�b�69��q#�θ�����&m. � 	��ڌ�%P;��}�ui�n�f}Q�Y.�bʀ�]�{B�Gdh1�?&�1��K��^H��/ŷ�h��X�0v7H���{�%<
��xm�V� �.xE.����.�r`,�<t��8�I�O�5�S�G����nA�+���t�:���0�c��I�xc$d�vď;X;��[�~����Ǳ����d�.Nﾘu_��I��o��J��G���L� �ì�sQ�Y�8��Xj9�g���y�}��8{��[ꛠÇ�����J8OTͽ�3Q]�Bro��6e��DN�		k��㠄��I�55g���7͂�e�B���j���ϛDs4º		�}728Y �G��������N��ه��~�H�b� </E���s�d�1&6�R��Cvw��!`�E��`�J�&���:��7(f�����ͬ�������<�1�W�q�7	'Ǭ���[=*E:X������8qa���	���9�*~�|/Ba����?���7'���6�@���	N�pi�2�Ce�h��bǆs=�(dq5�@f�/D���Z<n̓76�k���4���_uGĭ��c7�em�G=�i��ʋv��tx*�[��_�{DX�f����8V��(��J�6��+]5(m0�J;v��HR��h����]��˔��%q�m�V��̈́�l%(L��K�M�������+��F����-Q�)���|A	X�I��G���;�&��C h]�ve�����q�����`�قZݕR�n�\o"ø���R02U���$㕆ƻOY��֪H4
J��еCJ|)��&�U�DJёe�x�q���D��̷�9�
�{T�d�����~�~H��>G���=���R����x��qk�;���s�U⡆R��lOX�6�XW�$UJM�_jV{����/������C-�<�}�oM�u�u��j�4N��;���3��Mв��,gL1w]��@"�H�5�e�b�w�#.J���:�}���Pp��z@��I |���Y�A^�6p���LnW׬t9�\1,S�<��(*��^���OٟӄAzY<�s�m��=ַ'~=�Χ~�����,c��,�H�q���������נO�^O0.j�Y|Ev%�RvTڬ�3ڿ��xJa>�M��$=�T��کY�@ѓp�e�`{�3}u͡�Ǿ�iN4�G���U�z���4 ���N�Ŋ��عs4 b����T�8V�S,H�[��O��EMI�--nv��������Y�v��Qə�>�VO��)�����f��Z������^�������NQ럺I���WP�]qi��*��6�N�Sղ�ǡ (خ���=�s�P���V�,�Gp�ꏰV����� �wXi}�@]t���ϖ��B��/X��2s����TCYo��~֌\��7�+�@úx^XF����#(�{}� �î�Ȼ_�J�Au]�G�C 5H�a^m0�E@�5X�B�"{1{�
��;�� �9Yu����:m��)b�����Gs0�!s����on�;�C�ÉЄ�b0��;�(�c�����e�Ǒ��C\>D����o���� YX�"�5��W�G�y�Yf9#�:r�kT���,���I���_2Cʱ1�i�kD�v�u�_��~�3�`gR�?����+���(8�^@T��޿�-UNP��e2�R�.Y�u�]5+_ШS>4ؼ��LV/�ma�~��iZ"Y�A�8�U2��jOnt>e��=�xM�(��$���s��!���%�I�;�^>X^��{ܟ|.I>� ��������/P藕C>Mh9��(��Y�d.V���o�:q�1�@t�&��Y���~P��(%1��5�d����<��a;�y�3�e��7)�ڎ@	w��X)�;�u1c���H�c6�����B��Jr�����}0;�P���1�s�F$퓖�'�o����k�Aǧ�Y.v�M >�r?o�:�QZ_�V�Oz��U�е��J�4P9J��b�&tB��h�Y6:oCB���K�4/���4���u�6�;���tn�z�0�]��yYl��_�Zw��gU'T���M�$z���ѫZ�q%�"�"d�6k��dX�'@kN��1H�7Cɜ�.�T#Ɋ|;��-���ϻf�cf]����AL�^l2�&;~�*�*���|��H}��O���Lɰ�씧�m�M�M�|�*O���լIa�Ӣ���[�h	ر� ��v�	��0r��t��&�#O��'#0�-9�(9B�mܹ�DM�{L�2���@&��߂};���Cm&���̻�Ά<�"�S���Y�s[1u�7)�:l��gd�>����H�0
]9���HܒOf�D��������'�G�g���D	���N[�����	�#�;��.�r'~�Q�)�K���-*���y���|��'^����� ց*���n�h�~_wZ0�_W�*ձ띵��܈�U�wJk:$��I����/-�+o��2iF`3�p�j����W6��T����!�v޻C�
H|�h2��!��v�3��&sONg.;����ϗ�+���FJ&��30�2��'c��6�?��P�m�31��,���TϰK���k���c����3Uw�7 �U��Uk�ęd;x�q�D[���ʍ�$̪݀'��ԯ��$�j�<]c)yr�'P8
�%�ݷr��?��#�����q;�޾;[V�l6���B}��K�	�Sf���s��ZW�)��̬��!*P�O􉝸P4[D <�m:�"-*��=�YQ��a֭葷��/=#E�6�� ,�m�5q	�z��!�
��%Z��R���bR�WL�z���;�ʑ����͘����]E�!y�`x�P�u�2VQ�� K��+�*��h��56"��G�?��% s =���G��V�F"*��Cd@�>?�\�4Z������29�?������� �3�̳7E�l�-�<�a���D�R�"�d��潲�tJ������gl���f�:yְ}hj������Й-�5�<S�]��Q�v4T}���\�WR��d�r�C^���饉H��z.�<�70���s�V��V2a��cv0��<p���g'ŏ��W����4��v�Ҩ[��)� ƶc�wUv��zu6��T����@G,I��GhH�E���n�4��0�L�Y�x�)X���h	�=�1��8fغ����v��U���)*�0���;�ҕT�X"J��>:����&��o4kP�7Uz�NE$0=Z��E��0}u�J����`�<���$x�����m:Ʒ0��6�^�7���8��2E�N�aT4��5�_��{gZ	�8n	hl e|��ϸ�(�`�p_�������{N7��L����m3t�2K{���:���,Y��b[�)[��Hન����o�|���HP�(��㑬s���e>��GD��rt��#����B4�[�O8'%�N�%��+Q4������v�D���;�Ji�n�[Ml;����uw�\)�0�L-2��sfO�_���E�Kur�J��Ȗ��n��4%��rzP����zaP��D�=����Gl�I~����V�[�XQ�)r��[���f>��Mr��7��B=볋��a3ҭ�iz��ݬs��~_\rH�^�nf�?�I-��;�6�s����aȯ��5 �"�^\�i��YP�f�(1�e��	��������!J����<&�����D�����^�T�pI�SO�x�௼��^
q@Y
�����O���_C�TMvyCq��'_�d׾kՔ��mQ�z���)�>`�\em��Wl}���2�d4W����fb*�:�,N�mSC\��\}z���(����VS�'�Q64�Ǝ�$d��T и�Q�K�
�v�Z��+��6�`˕T��i�����s�
�i�1-L��q�?B����*<bb��@��jf�.���v�#T�VmU=|>"V�U*�&x3_�a�4�}�?�Z�����=gTq��2,~n�䕓Q���Y;4ϠA������٬7�j��Y���J𓨘�yt��� F}R'���<�G-����O��!��r����ձ=j���,����0��;P�:��jރ�sJ�]MA�V5Q�x~n4���s:���}��.���P���=�U/��H�k�{��9�v��=�l�-�P�+_�*��t�����Ȁ�t±/����ڶ��:|�4`q|�K�,�JD�&జ�y�R��b!觘m���q�䛼�y )��)������qCf�w
��|d�`n�n7�l���V��O����ͽԺK�C*���f �u��|�CF�e�Z��������+������>�u*�{)�� ����.��wi����q�Pz����?l�)�my��=#�Z��@�Њ�:<_РP�~]����D���l~��Cdvg�����/V�=ں)�W���������PFl�~��S3�bW�c_��KA��#v>6V@Z6��s�	�����hg��oOk(�Z�>��p�<e��]�6��������ٗ��b�G,H�.�퉘��5��g�}Z�K�y�����b����=�1\!���.��¤bw���3�<�`,!�l5�I$Ґ����2Ql��Sy��k=���(�wP�~��ma ���G!ѷ(�^-���K��5�'a�
G4;� ːJ�-8�zK�ֺ��Տ&�[� 1!szܟH�qv��3}�3aڳ�e+=��۬��s�R�W��'��x�H�ѷ��b%�]��<�E���V'���c	��u�mG�ߙ�����E��`:���I�h����3�7-�e�>�{El����[.Fwh���x;D9�<��	�/ �顾���Lhs�j�Y	3޳� qa%�+'z���W\�n�%�lIn;�{O�%>�<g�?�́:َ�{�7{�Z�q�/.��Z7hW.Zd���c'�B��ܓ����e�hW�Y�-L��v]+�ne������s�u"?ƈt�)�� "���
��B+q�����z�S�$$�"Hʾ�K�2�������}�����z��.����yV�/R~��v�m��v�;�k��E�Ji�ځwl�kL0�0Ƣx�'[�\�G�&�Ngmާ��7ܐ.���	5<t�(��l�������?�[�4x�����1H@��Y�فGx�RÒr��Ezk:���}�c��hZc�4+L����4S�`K6���`��HXʣiIX�?}��򫫌�m����nWꜘ���dNn�x[IOZ+`yN=��>1�jTK��k��m	%�f\S��P�����e>^��Y��/¿����D?��'��4��\�Q��~��ϳ�j��p29`��Co�>�L�3��*5�}�Z�E��bm��M����D�)�5 ��Q�>� ��Ĥ4�>	��;h=4*4���i�ʅbs?���kt4G��f2Cޚ�a��N�o("��U�h\MT��&���cQ����s'���@����#>��z1�XK����^�[Mj��.~����c0+�k:0j��(�{�}����JɊ�����/1&O���vO=�r��I���5�����ZKC�ԸeU���PRh�� 6R��L+���-&Tm�f%%�6R�Ŀ:I9�xG��ꂸ[Yý(S�6�\87c>�A�)^J�6 �~6�D�X�.��)��!����z������|��)� �"��u��)�Pva�tY�U��v��@�&b� 0�N�s�XĎ�x�ce�;8�'��x^�r���s�.Y��W�oO�B�:�$\���u1�wTn9ڏ���eK�#�G�w*��ڜ9�.d@w뒪���c.O<�i��+~�����Ztq6��Bw1ʖ�Gk�8 ��Y�����N��>MJ�k+�8��6n<����`�I�$�5t�o���>�
M�V�����85V�LT��Dh�uK�[9鐵���Ơ�W�����.oWo���  ���6�=��:��7rRC�NK9p�_���Y�����7�r=��S���rʑ�ya�@��c������ hS0��?@5�v2�n��3rZ0��8�,t�Jb�r���ٿ�wr~��?}9�ը�;�ԍ�����S��5���5�g�4��*C&Z\!U���}xXqP$�Lr�]�a.�B���hy5�[�bl筹՘��wu�~7��qL�rR�E�?Ƞ��k�:�R��W����UQ"������x��q]�,I2�7F�<�7���kC����DH���l�wH��`�Hu���O�ͫ��a�O���k��B�_��x�Lq;��L/wK��KL)��r�N�� �R��r�݅�Q<-��p�J���C�N���ڦn����fH�T�gsG5ϥI�Љ+�k�Q�8�����Q�������ז�;"@�"Z԰�4΢3�K��^�Lr��lE��Rˤ�"���8�)�\}��՝tțYh#4$)�81B/�4���݄��ԇI}�0ML��x˛�PF$��%�!�6L�\n%��]�k IG �s��8��A��
`Z:I<��^��z���uzx�g�bղ8�*���uK�otS�l���8]۵Ɉ�!�22�kg]�F�p�e�.����"g�MY�e�
��T����h���^\�U<d7����0�.�zS.M��M@oT�s:)M��:6E��Mw��y$�Q�O��M<2�g�ޞ�I������m���v�������t�>:w�=���`���%�G]��������N4X����YŻx�fT*�$����^Bȶ`D�Zyg���tݞ1�~��vy	�ͅ��n{�����R�5����T��s���r5�]�Q�0���a�ǹ��/�$�ADV8�D,�q.�����0>�� e���ҿ"��?�ⅎýݪ�f�� k8B�@�$ܽ�p�L$|XS��]�,�hrx��-~�m_�u�����aWp�݌?tm�?����>�N�|�(�%�섺��L%{��[��Ɯ����s�e�_S|��l>`���fM�管��Rvo��h���嬩�΋*u{&��̔�zI����ǈ&f��aL�8�z���Gy�}
G����U��ׇ����o�EF���Y��F]o8�i�_��+��O��J_u/��P9��T�\ksG�m��5�N|�ބ<<J'A����\TC��"*F,lg�F��ȩF��L.2�$1e_�Me]v���	�'���>`x�EFhҶ�����x��4���G,�Љ ��G��Ҟ��>�a[ȶ�	��0c32[Ӽ"v�8(3��p��|��P��c���7�[�!��^�x��Jup��L^�
�����'�ެ����#��K�ԋ���+�6���y����!v�A���r����ʯ%f=.�؏��#m	H�nUU�)'!�v"�#�-����b��Ư7�zV@��LQP8�����E���9�F��u�,����g�t�4��3�*MWoH(z��a/�z�'_���تS5Mq�'FИɣo~RE��ܒH! 6�j�#��B�#��y�&�L͔��q/��~eMq\f���9~��ZyW$%A'�����8���#d2�n�;Y�����ZSMڴY�C�Y�J�q,g,כ��v#��)u��E"�
�/>�D���½���ZTR���&`��=K�E���Ў�2��XjB�f�2�u�H��a��mj�p���?�
����]�#E�]�n�W�\��	����0a&$��ɿ( ���ݙ�9�{�4O���S�^"i�oD?2���=����I
��0�.v�T�ت� 	'�vZ�p$}��1A�����F�a
���в
�i�9�$��Nr}�Ț�qOUvլ��P���dG迠�\��D����c�&��2�EHq~�3䉢�k���!hv����4���������n_8nn�ȝ��.� e'��C����0�a���fܻ?�I�t��w��Լ��#���6��:]DT��J��+����TT��dh��o"l~��1�w5/z���c�U�WdG��f��퍍����^/�l�[�'2ʻ}H���<���T<�uŐ\��
���$}��QI�=��	�E9���z���8�d���?��$[����J�jzW;B��ޙP:&�y�S�ey5���%<XBB�'b�"oʹb��J5_ :�^��� ?[bL�p|��]u�A�dk`(���R�ƬI�ŧR��"RqS�O�� 	
��".��A��V4L�@'��]��a��,,Ž;=t \4��:����\L����G8������(�xgϱ&}U-�d,0���U��c_#��ȗ�H�|���N�O ����e�y)�h�rc>Ȕ���8G[��<"�x����8�U�_'�	<.�˻�_����Ro��7om,�*|]Ή+�XW��p�$T~��~V�!������?��~��]e1њt;t�@��e�R����ޭ
EtEz�4Dz�rX�G9�����~��dwXj�(U0�T(J�%�2 #q�X�=C��qY�� �&Dm�	�72���}i-��&�����e�Pd��O��+�z9��%��ビ0<�ƀ�a�qQ!ɟ����k!�<�;��
�f�-].�)�x�ȩ�d���xd��z���� Ƴ�|��[�vl^B+Q�J~# oiJ��d��Y�7W�IY�3��I+E24�]�"v�7�� I�gRM�zg`�6�l�c��Ke���p�]��<��lUݾ�e�N��%���Vl`'D�֜~4����7�=�3K�Q�W��t���}���˭G�/껤Bx��7V�&O4��|����"���Bm�i �=�_5��g���ڂD8�1ץ������`oH�r>9�0?9%���U�0�G��em� ��0[���I������&��p��v������L�'�����\������s�i��5��ĖS���X2��fy��ز:���K��!�v��塆�#J��ae��N5���d�'x��� �ָkbb��_��I�w��gN`�eM���*x����r������P+�O��k��fw1���5=@��r�[�at���>���w�I�V���KO�&����0�P����.AX=j��� \Vv�g � R?��������@]��!8E��3u؇K�}[�k��Ҏ�ya�����\2��T����/@���O���jZ���O���L�&F�rW�ǔ,�Z?O�B�aw�&p�iRV��.��ǻY�=G0S�v���+���Wʞ�[��2��5��{�TW~��d1K�^/ӊ�P�D�RO[Z��$����v�e޸���Tay���@�P��i=�.�O��:*�q�2��*��	8!׆q����K�+Ϩ$�t�Z;���a���g�{/ 8��i>��5�d��+v~�g3����E�¢�R]��i+��VHb�c�u�&yy�� C�:�):#%]Â��bx	�j�-L���}�H�i�.�}�\;H{ɜ�FD¹��8W�r���0�}G�����s}�#d��-�be�?}�� s94{��rnW9Y��c���lC�k��es�쭒0q��+9��O���νe[�Vmb�p3e!m���Q����n��o�dK���3�=���:r��-���;���
��6%�iKXey�CV�����tŲX���棈�㩧�.^E��&�*�����^"�ˌ�?�iҗ��W$~�oj|��cBǯi'�������J��U�y��qF��h.��}���5 c����b�.��u ��1'�;�p�nw T�� ��o�V�nI��Zd2�~f-n�&��X��ec������CL�_��u[���؛ؖ�Y�P��'�d[�c�w���T�>��mZ?f���­�e�WO�� �����s��]=q�0sW�{2擼L��j�"��	PII��Q�cNԬ��+�G��zÄ��T;4Gq�n�����<��;L������6q�!	��l(�^��R� ���"Y7�v����7z��r�V)F��'��e����͗IA�e�����1y��Ce8
�暱����|I:A��Q�K�;@w���~=t�Q�;/�3%�PL�lX�,��{ey��y�J�z\7&J��!@/��Mfי�����B�\�1#�nÇ�)�i��$O'�������� ���~��͓�i�'�i%6V,�_1m��٨]�k�X�' ��k�"#fr�5��^��-NG؄'p�R"r��y
O�[JS���$���[�q�t�K
&h���
ψ	����5
3��{qM�	6���sK���*4W�gx*M�#�#�����X���z��.���#&����UƆ N��ߕ�s�S�Q�4�t��-�-;�T�w�`��@mȌ�<v:�Q�گwG&nO�����>T��l���%!B��iЄ9�x��p�uͤ,Ӏ���rYYV��c}b`uJd �y/��7�J�Y���/��;�5$J�����44Ы+F���<Z�PS��J0�B[D5����kx7�{t�Ш�G���*_nx��-Hw��l�Ep
��*'�!�d� ��������\��x�Zު��1�XH��̔#���[.���i3G�A՘������4h��M�H�:,��|ڿ�M�q�'�}�P*���$�5%=�n��٧�G��\t����	?-e���*|PS����Tٔ��Y�-�D"��Vs$�N,np�%�F-���^Y~A�J�Z-qķ2�E�j��E���.��������B<�$C�
{���#��{s��R��y����s�&�˹�Aꯀ9�4��ydCԀ��3W��c�^-�͖h���0|Ovs��!�vn�ZV��,p:c���	���i��੶�d��6YV�v�"�y�F7'�8���cI�~��u�Q3���J(�9��g���Z���V8��2Hd�L������NG���@�x�����֝Ma��vD[�	�U�w>�K�ill��uw�k&��Ů��E�)�f#���p3~W&���X*�m�i0����ߗC[.0�i�B���ɝAM`5b�L����*]�'��2=�ˌ&'ɝ�|1SϷB�b�p�>�r>M��O�����H�B�q�^��E��t9_�� 3M/�X�}� c�98�����:�N��:e<\-�Pe��5M�iՠ��[�8�����R��?�W$��G
	��8Y*�n�Ip'�������,-ѝ����ؚ�e.��»s1�}Md�%K�:^'�q�c��0�ǖ�:g�Ҍ�|ZdP�����_c������M�5��l��`U�r�[	,�|!+.��oQM�_���U�DCoݽR$�A�}�iݽG����8�6��,�#N( oZ�ƠmE}� ����l�Qv%c�Z<�fheO�f~�/��}oV���E-T���}4��9I��a!󣀺�A�	%��Ҍ�@Z� *M3#����\.$t�ެ�X������t<����Zv���?8*'�?= U�<����Eボr���G��$�M��FЈ�d���I��<�����xT$�Bz��q
� �]B�Wz�+
��r���~bp��.�pB��o�ٚ��.�M^�^"�!��"��G��z��^���S'��o�N��ٕVB�r
��1,b�$P��8M~;���M��p�1������<�}a�� ґMw��-or���y�����i�`e����]����>/oB�M��}#ȉ����ܗ!L�6�m�b���xl�D|]�U�8��������s�.�Iv�L2�4 5�Kn��$�����Ʋ��C����5[x�.M�@3��& V{�*	�/����;h��?�%��. �pa��h�lJX/;����^a����րeF�E��j��C`����ԙ�l��I@��%h[�l�?�}=�@>�Ð�n�l�^	�it�7�(ܖ���C'Rr_�)���MXrpT�&}�zr�Y��a��nrB\QJ{����k��w�xO�HQ�m���fd*B��BN='8����I���K��P������YN�ӄP��JV�1�?�:a��L˭��Lw�����k�e�U`s��t�Z\��U�����C,�=�����k\@c|�6�Q<Y��Ά�VhCp*|��g�����h-��,[��@ �w�eA��5A��x�� O�1d�$8J�%`���|Ji�����=3��q\R���(�]��rn�l�@��l�����oh�����]&�O@awܬ|��A�R;JZN��h+��M�W���k�5E�K�zx�4�����&�Yp*�hiC���]͙ԑo�2���"4�~V�֒# I,�t|��jk�s�kh�1h�=�Ы�޲�Ϡ�����v�����*Y��(�v���Bzi�@4��Kg�b�缺��4vG���i�����cI�;;�Q���_>�ѣ>���]K�_{��RX�)�xƭ����C,���#�e����6�����_��󜴏�5þ$R��Mn�)��]�@Ѳ����U���_y�t���G��bc������:�N��D�dP��C;�*�Bّ��$G��,��IV��B�G�\o�ir�-Cr��Ѓ6����Œ�K�ob"��/y����t0��2U�^�)I�M�kdSs�/s6H+�q�[pDp�oւ���#يu��߆"��c]s&އ��O���+�����5��PI��d�8/�֜ڕr��.�{�i���,Zr��R���Ѐ(��`3�e��C����͋�b鼪�=�h�5yu�If8����>  ���������)F�#�^	��(�����;���Ln8����g_�_�R�� ��|��]h�JH&@���Gf0t8Aî�7܋A.wi��<�dS�oӤ��i����3�P	�K"�{�n� �7|*��&��p e8��}l~���TE*�tR�>����9�Y��ȚoW��)e_e��}��>]ʹ@ea���?�P��K+��w�ㅀ].*�t���7އ�@�"�o�bd��q�U��{�k�s"�H�z��L��*]���}��Se~��-a�c�MB{�u�AO�c��t˾�x/�3~<����F�z�UJ��*&-f�������x����>��.�I�3��@� +��ݺߘu�Os�u;��QO�6u{"�c�?���*����ZY;�󗑱���$��&"�w]pP՝��_ej���-A�I ����g?H�Ìf��=UF�9�1s_� 6BbS$1�3/�����Pr�~z�Jr/�Iv-m��E�&�!����ZMi�W�C�J��juPr@�2�jԂV0�� �Z��,��X�yL̬s��	��m�7���+��Ӹ����L�E��Ŧ�س�>��u�D�Hqebn̶
W�9�g&(�6�^k &$����ANS�xm�u��g�-��l��9c~��#D�$�7�GV�Q�H��5ir����
�>�4m�����Hg%>��)����U#� s��́^��M>Ϭ�!��u��'TM�k��pNzh��_,�{E����op����������s�	�IX2^��{7S��:C!�O��қ��n��g\"yX���C�z�׏,˞��{��0Y���?|%�E��^�=\_���s����/�l��2 Ί~�T���A�.`�z~j�}����R�r�pxK���;�U˾�ݩ[�N�n-1�V���Րu��":#j��X��i	�	h���B,�tI�\[\�81�Tb�[~���9i�a�.UN�Ź�������"~�����p��jD�ߓ�AȄ�P8ڰ���1]��d:
Yj\�2Ʃ�;c�z��D���B��ldR�?�^��-zؘ�=��g�5&p�׾��=���\�U�3�6㣔 �"ZO�)�T�M�������X�H����%>~ʉ~�KX��(��������u�sB��Oc�E�O��H�5�u�_
������ty_�u~IX��8�Н��$Q��5a���4�6x�f��zmg]H��Yl���T�YbQR�Ğ��8da����ˠ�L\��GEx���¯����Ac�� �;^�>��L2T�g��F@��\�z+�t$ �¯���ɡP|.��>��	��kLQt*�(�g�F��� �M3�LM_�n�3�+P|^ف �%�W�?Us.�����l���F��r�zw.���Gfy&����i�T����1a|.iTvo_-4�-#s�w-/$�%���
�uK�(�6@JY��5�-���gD�p��3AA��h!�,8ڰ����"�^��4�$�x�<Gu�u�"6��˒����Z(�N��#O�|]mop�G)��O�� ���)�c}�Q��j�gP�XD��=���8�5��!��hy�o�1(��S8����C�����<Bm�TÒ��ˌ��Ԫ�]�8۶��z��@B�V�9<�)�Nþ¦M~�-?�GT�g!e5��Lh!�,k�U*�^������R��w�����ZSg���t7<~�DԱ�!g���6�M��2c"�o���6`B��O�Ԁ]�P2���`��][P��[�l�4�y��Ȑ7m@M�M�|4>�M�+~W�h��^φQ~�A�{�v��؇�k<�F
�I!�i̝/>آ��e��:2���r75���w�Dcؕm��niUr��S��ʟ˸H��Α�������FQ�/߅!'nZ�q�XX��5��~�� �b�%~�O��&�*_<��|�?�D��L��I5���w%�0s��Ps��ud"/_�712���MC.$�����ה��N�7m��pؤz����Ƣإ8 � ����V̻��0h
�ұ��z�c��d�j����:�H�79ۨ������O����l�������Hx��9�}Fe��b��ԑ_"7xf��d.����`�W7�!��ð���o��t�|�`USXn�GJ�+�����_�G6���݂����A�\>+r9�3�;f��*�$�ܤ
:�5��YѬ��*}X~�x���!{���N�4o_~˴1gi���ȡ�ͬ�͕�mc�\
!TIC���
͉=�T��iy~f�u<��G#���<Н��m,���)e�Qk�]�O�L�~N�-���^z>_�(��	8����b2ͩ?�j��������7���`��wE��D��z�u~sMT�@v�;{?�GW�c�CM����E�d�@�?��$e�i8Gx.aM�gڴa���]�G@�{{Tɏ�ܖؑorFZ�{�����%��{��y���8sHtr�X�:������1�|٨�1dג�����r�����h��J~=2ȇ�j4�J,�ea��݅
qwL07����K	j���۞"��m~�`¹1'��u *B��&�-S�c6�A�~w4M?��n��Zzl��M�fu{�_6�
xƎ���>��
��q�yM��a8棴���E2e���q�"`4����}6֡��Ț�D��p.��$�����/�-���#q!���v*|0wtx��ol�3���C�USWr���0��m�\K�] ��3���|��P_�	KF!��e��_(Ґ��#��xcR[�mPog O��� ���񠎚Ma�|�$��h~*(}wR~��
���~B��?	g�	��8���k;���(`��a�}JBhr�����*�+�l[��'haQ@�����tF��̞[�+��0�pB�(�A�>�)�J��sI4�v�L�j�>q��7��u.N��!�27�jD�㳿'̟�+�*��e�%���e����q�-Ը��La++=�.�\��|��t$b�uC�{��3U`b]2LW��wn'�@�4�ʯ��9��ެO�u����L����S-�<ɯ��NV�Fo5��A16m�V�	}޿�%O��I�W?����ȏ\� Zz��.���5Q���E�7�R����� >�|�>M#�����-�p:9D`qx�%�G\����>uZ�/�0i����1|�}v�J��&Ћ����ӳΊ_(�#���W�+:q��I6�͊�U�c{)s\������E���\��g-�Y��;�k�_f���Ezz���B�T˵Vt�'\�9�$���q�"�����q9��l��;K�� 1xn��>�e[�E�C���`�a� }�$��	�Y�g��������d�~G�?+H'�������[f����P�µֵ3&����ڙ�e �6&�L��Q����'�q��	 Z��R�s��ϯ�fE�;�n�M0z|�<=���"�R���x�h_����mo���qbX����q~���>�/�z�oZ#��Տ$`��+�`�+�
}���#7\��қ�\�	�A�v�N��Q���Wx�D���'��I����Ko+E�e���8��jDE�c��Ȟ�S*��[ʔ��c�q�-tz�|�ns�
�����/@2�6�`����%���$Tf�����L,�h��_�ɩ����7�<(ɋa�����[���1�)��_j��?
��+1��J�m��$�/��8�@$�ȥ=/�֨,4'Ŋ�Dc�wB�!A�۝�*���8\���9�.�b
�uoZ6��W�18a��Ole|}�.��W�|5��i,V�P�5�������gTZc���ߎ�����i��h�v��.3�ި���}�`FF�}�ϲkN�?��Q��U��a�����0��'7w�MS0�y�v����>hҵ��@��X�4�r���H�w����iV�����!c/�*��Hu阫�a�:�2v
�T�d���d�vm��I�9X�d`[���z~����z��F �I�����̓�
�
��8)�82H�M}b��M��zO� �J3���dj��YQޛ��zs)
��6��M3͍A><��o��ۡ�yJ��/�-�~��]�n�bJ��w�P=�w>o�`#�k��y*Ց��[�V��yw?�#g�����t�	�+�f\���2���>�˱2YC��0ݳ("MXn�W��Q������z�aW��o�x*}�Nw�M��O&��n�R�L�RxCm��k�NT�s-��o���ق
�+��Ǖn(��g[�����L��/]ْ]+��������b�h�sUҲ�d�3 �bJ��xf�1,�JH��sY"."�#���P�,mWT�<A��auj�°�q��3*��v���Ho�f�\��]B06���KPt��/�2��. ����D�p�j�,?ԎR��R4�Ԍ����O�CO���	��"���YS�B�]v�i=����=8@L-
ۘ4�s>�}������g�ex6�m2Y$�O���h5���h6]�9���;�X���T����P�c�Kjĕ��>BW���3�Ȑ y�WP�O?�ԥN��~����� ���jUh�lNK��D��.���g��34�T�����>�{f��/��H>�e&E~���q����v����[X �/���{ڑ%/�p�L:I�j���v���q�>�2Q�l���L8��e���^�c�a6����Q�N�O��&�Н�/��#���%N{�T+1�@���2���.yje��ib[�?V#���FW�Zf��=(*ژ�_j�&��}��pK�o&���2w�r�QҪ��*��&{�\�ȏ��.�B$�f�7�K�嗗}sd��-�̰��RȒ�!:F�k��u>���2�Z����6��h�dp���m�y�8���EU��} ��3����1��.������5�8�UM�#:l��s.%�#�`.��~r��5��jV$J�@+VݜX��J P�\��0�fg��#�u����� ��\��"&ioG����,!ɨ�q�\Ձ���d����x�خz�y��^*�{�\�כ<]�O��9f|��?��7�k*��Q���!�&Y,vJo�}gM^V��,�	���n�����j�$�\���$���9�WA�7�$������q���Xĥ���k����]Rh�(�"'�o�W��=N�ʡ���;��,<�!�{�R��4��8UD�L_��X�N��;Tl1�W,.�CQ����6f?Po�@i0�}k>w�2qS���[ܧ�]�8&����!��2 ���q��� 1W����B�Ce��A��I��� ��Ӿ����#!�I]b��҈��^Ă�w
���"|�,�?*P>��i������~������ex�a莸�?�w�$b^���}�i�ȝE��)���MԦ�[��seV��g���Qm''��zL]V ۷u=%�vf�u[\��{��q�d,8ؿm�������Ȕu���@M��Q�`ߒס5�I޶�.����*�;�/�-S��tu.|M�L���;��'�PŌ�uyg<��1������`F��u�Ф����<g;�ܤy>t�}���Te��H,����LR�����CY���_�Y<[�{�6�un�U����i01��[�<H5}�d��N	@�x��PmFͤ�7���W�[�|
�i�8�v�	\�tr���oއLp�����&�h��, ��\>0�䠡>RV��=���P����<�.-�0��l������p��ӕ� ��#1����z`��&+y���ڬ~9�7���u�B��oM��h�~5�#xfT�Ό�t�$RJ�t���*���je�B#1J��v���=���0�Я[q`�}6���[���ؓ�
d�E�(��5�`��l��e�3�Ay���A{�+��`�6��Bߌ�q+�ٓW���m��:��Ia��I:��<RSY���#q<���h����t�E���$3,>l�N
�s8z�r��gE6�K7/�����˞��̬����`��wc�)�t�I�q�}�y}��gN	n����Q��d|��%�[��|Tu����]�\Gb�N�XyQ���&��\8Ŏ
/>���������5)�[��o����e�ӻ��ʝB��z׼��¿M��y;EO���Î]�B��:�a-E
��|�0eJ�$��ǈ���u�UʭE��K�y�-��휯#�@�Z".���	qC�=g��G#g��Ÿ�ZPL����2�
|��\��뼯̀����ŃY���*
%G��)��0�.�4�3�����%
?�	�E,3�ߜ|�Qb��:x��ύY����C�^|@��ɘ�7y�ҷB��8վ��_�d���03�`�k���ŭ{��s�������D�"����:1wƖţ�	
���ʎ�9�p�O;��I��H��:���'�b��7� ��-V��[؀EE�u`u5e�w�i�SҼ.�-� �5�w���c������@�����������>;���A�f4����$�)�O����؎W�GP�I�l��%�����}	@_7�_ �gK����������|���Pʉ��O[be���UL�a���7�Vp�R�M� ��aq����e؁����4��&�P
�ʇN�$R,�XA��.�'y��7��;���5o>�a���Ղ�e�L����D�2z��|`{��{�+��>�%����_9<Ro�1��~9.��d�2����D�ii�ɹ��a>���W������bc��L�*�7�s��Y ��<b�ح���,�r��d���[��a���1�`�׶~khhm6�J��D�qiR���	�a��uA����]3��)���1N�~-� �>�>�d(RR��2� ����L3;����z@�Ҟ��ų�B��fb�e�q6�}W�i8C�l�ib������E��uB��5C�c�CJV%Pm��q�Uq�ڝ��$�W�N��ǂ�U�k���Y��������C�'����6�u{�>�K/2?&����'��3�/uȿ��Z�ǟ��!h�b�)��9MD'MY�A.�K~��%j���h9=�~�AjȳWG���[��VRB���n�?���\�ƨ���&o�d�چ��? �&�#I~��ԑ����J�`�y�'��ز.�G�g�T�e�w5n��u��"f91o�%9_B�����QV�Չ�7U`�0\R�V�c�oL�=#l��}"X�Be]�,���w���7i֌b :4�
S����d�7M�lL춯��#���˃A�@i��R�tj W��A�1-w i�ld�뻝J�ə��)r%�5I�)#A�{�%8��)I$���SO`����Yv�dT�%6���A��z��L�y LQ��� �ߔՏ���J\�G���E�}ty�`���8����r�y�L���G����$�t�?�tlޥ�-��y@��˪)�*8s���0�����kL���B��R�ݒ����U{�@]�8�N~R�+��Da�nk�|~Bח�<b��9.V�a��:s�޴H	�����I:�����ϼ�{OR8��k�5t](1�|�"p������.w"U u��
Vk��B���ݪ�](PwT�ԯ�
X4f�|h�,��(�մ���^������%k@�#=�&�0�u�D"��m���ҫ�o~���"ҵQ���T�qΙ�?mP�X�S�]�gU_��|�c��{"w��[�3������XA�k>'�
FOP��X�b�O!� qh�/���u�@2M��w�1��0&��L�dJ��!V�5a�j�Q�CwB#R���r;mv�}0n*(� <,a^���N����}1�	����f�JS2�o?Wz�\Qw7W�)���h2�}�<9�c�U~�c��@��}	��� �9E�zc:U��J���c�<��L(G;�Υ�k�ӂ���C)5��S�j>��z]����U�Р�¿�� ,����ڙ4��j���=����j�M���P7�J����'����>����T��n������~�s�`L�[z�����4(n�����}��
ڭ	�����En�J��χ KY���=4*}j������*c>����0�iD����k4`�˦��a�f@<�i3�v�R�g���{��pe���])+tc�ɚ����b䌘ahɾ]�*�T�p�?����Ȉ�Q��{�C�b��иa��^Gu)Vt,��53�IIݕ|t�g��G����5VЬ>��y�F�ZZLF�H���F���*J�d�Y��t���ɂ��*�d���ۂ ��F������V��E8����������<��.z,g�R�q�⏖�_\�KEU�,7���X��P\>m��W	/Y��'��O��LI�a�ag��4b�B��l'ѳ+;l^��3-]f���&�3LA�,��a$!��!rp}8&�$�|@���BH�!�����J\Z^B7��u(!�	�����R�Vβ�ڧ,�,����r��8<,��Qgu����,t#��9�U�[n��]_s���X��{ (2��K>���ѫ�j�����i���ĸ�'rS�h�p���s��R�gr��0|l��[DR�
N�6��F6+v��К�u
�F�O�'e��*%ы��lE狀]��ύ_MJ}�L�&h����P��6�H�pbPP�x,�Vr�P��*x�����4�^����.�mG*R�D�>���p����EϖX�h���5NǴUĠ�bM�ju"�Ƽˉ��Io��@�?7�0%�u����:�s$|��ᘥ	*җ>��o]����J[t���K�3�w����|>,��I�}�J��Ě��XB�﵏���Wmz�G#.=���C�qw�.�,^�u�G�4��R��Q����n���雏A̦��GZj�i�"v��P�2�F,���*i�ܤ^K���ț$	=��}�4+4�i����<���}��
�8�i-u�3�?ձ�MR_ӭ���[f�s�	�:����Aq�Ӛ��B��n�� ���f�.�Om'Ǌ��m~���Hrm4 �O���0`��A#[��C�⠖1H�Q\z��ʰ�!w0�.���Sd�T����a�À�Cf̄�������9��>G:CF*���*��
6��jȀ��!�ޠ�����C�*�}/I(U#+$�'����O�&�I*�a����NƱFض�'�Oy�Lv=B�����,	S����pJ�.�>�a8~�2�v��&�<U����[�^637�mT=�a��]��4�:.�ǁ����X��¥��y�i��3��Ɇsc���}!G� ��޷j(,�H���5���;��6�8~�$��ϭ�7�`�|�'^�߱;�D���l�N�x�:pf|z}��:��6i��!!��f�����^�:\��,\���Z�(3^�}�����A:ot�rt�,��/�x�,mV�.�jK�_�6q}��Dc�U,^�N �Z!	�N��{�{֗�G��UҸVyُ���.�D�*B�@��"��GdWj�O�97��<���Q�[7kg#P*�(^��l�?}�����Q��&����d1[T��(L,ƅ�~_ov�̤����Z��p��)2��q����&��M2W2��]�(�*Z �&�Iy�Y��mgG��٬���E<%(Ȯd�g;z�(�ʥaa,��2FMs[�-��ޛE�qD��.<��x����/b�$+�� ˼�He�����T$s.��c9,��3*Vq:Z��]�X�;Z$
�.��L"��-���O�/�n�7^d�s�z;�;ᏺR�!nZ��Ǥ{���k��0Kue�r��5�ۚ��߼����v-ඖ4�<Oao�Ʈd�\�C@@mH�,$Z�)�������aI��-��6�o ��ݩ��e��%���"׷>�Ӡ$�`��; H�me����9xH�����S^��6'�n����l����x�%�6�wGE+Lf�#j�(9)@])�ţ{3\�̫
�w���#����gK!lr�A�m�|\]�}!"d�@q��SU%0�*@�a�g{��}�����2�(�� ީ
a�4d�dE�7�v���?+[{�d\^T�8��o�zm���eW�����W���0q�ŏC������K ��c���h�O96=�V�b��ˋ���)�e�!Hbap��7_�${�G��K��|�/)��Y��TYt�n�^��>.��y&/a���f��-�FUJV��Ŷ�27������V��Fuq�OA�Kcq���;6�eB]:w]."(5��PB{�Lm%ȃT��^(���zSz���@^ƌ���_�W2K��6I�����	Q��L�u�.��4NonǪ���(����/�j/�tx;,4`t7OY�x}�#6o���� �ؼ�a��t��$�
�I���V\�`�]ۂ�V5D��X��#\m�0��{��_K#f�_v��b'�F�Z�V�ML�>LC�&�6	S�����q����?hY �Q)�4m&��k@zMEr	M[}��`���G���K:���ՃlPY���!�P&�h{���n)j�l�sTؤ3�ڲ1&��n;N�F�q`'?�p$��2Q�|����m�߯��K�d��W��f���0ϑ���^8�q:3��ьȵ�&���1l�7��xa��ս��`L)��x��-?�1l{v8h�0���6��R��n��,-0)W�[Ju��F`E�}Ë����b����FZ�k Ó�̃���XF*�����k�FI��\�#�c��?T����.��̙�-��*N 25"�Ѷd�ƍ���>nP��"����̨�O'�by���l.�� e��b��^�kI=�2�{�ؒw  ���>�o*����q����k��Ζ?p��B��=FJ��F�X�`x�(�^^A�F������Ͱh.Bk6NA)�h��Q��l���z���SC=߉r3+�i�`n;���	�V��8A]���lWM9^�T���'镞l��S{�V1�������D�լT���pa����e��c2�_�T�j��zB�!�K=vQ}ʈ��[�����%�z�_O��	�;-�]���Rr�MQ4-��h�o01�>~��+5n��U)��Wk�B������x����:�,�p?�!Lkح߉��/��g_������7�ff8���ߵ��w+�C���c��҆��� [ġ7���	5fSu\���b�)�܏T������Z\DtiwZ��r��t�8����p�ٛ�=�K�-~Y�ݡ�2��=h��唳��i!ǳ�wv(��"P�!?c�o>
�ڙ�h={V��'��$�
8Wy�L��t�cn:���p���Tr_�1�=ĵ�����r���Wez3����|^�FDP;�Y���f�sC$�x��'�f�U=���c�_��A�Bh�}�c(8O�6�����GC�����(;�9q�~�$;����]���!i*>�9AC�P�����RRRT�BN���DF@ �xU�ga��E�����T�CŴ�xL+ѱG����E�1|ޑA̆T��J/��(09���/�w��w��	��5 '�N��R��bW��^�7 êGj�.�QH�"�x�V��C!Rk�B������5B�OB�!(��a��Q���8d�\8�pA�]���=c���������q&��i��#(��o,uG���ē�OݐR"�YZJ&�#������N�jэphT�3����3R�¨"�_�>i�[%��}$��!��{V�0H`����h0�S�ѼO���j��jY��|3��!%�;����"�ݻ�}8�>�_��zL�W/������bdr\u�Tjlx�c�V�+�u��*�ai(Eپ�+�_G��Qyi�=�ϸ/�x�M���ݷ�+���MHt���o��H�z��栥d��oj�*.s�ÿ�n�����ߐQ#8^Q����O�N���y~���a����7�q�R�,�:,7^=N�C=͇��6tQt���+���6��?'[�pW��!G�������u��#ˏSS�t��r�Xٙ�jq2)�!�DN�(�x����t�u��Jj�:|�l�iG�Xxz�8�b��7�_(�S.8V�{@FE���\3EB;���P��I<�(Z��[��b>���s�L�+�)H�A��D$d��oT�A�^+],�}H��m��~Z������yYT�uW�.��X:0CX��P�j�Yy�`e���IН�P���8}N"{)+#ғK�I,�ݣPPS�Uʑ=�"P��o�8���;%��q`A��ћ��������9K��a�I�x��b7Y4�b3�MP�*Xg�I����vM=�Xx?����?����է�ȸ��d�C�ߒV���҄*�rՆ��CU���R��gh� �	��X&8`��AT�cM�fg� �^$,$Pn�
J�=��rV�+,�F��a���6C��% �C�(������U3!&��]G������$��(`��������w��(�A, �k����'��Z�9�c�ݍa�z�I��*7U]ܶ���/4��sKKL?q�O���Mr�o�o;�h�<�U�a�o4Iw��3���*pQn��nh���`�*��KD�dZ�e�����(NK�m� �F�GI�`�YRm��G�I��>lJ��r����'˿��M��1����aP�6��!A�X�<��S(�{W�����#�����v��� �Ϥ�v�؁�A�/�d}mbؙv�"��G�l�:���O�Sx�1Ș��|�4��o�����&�.	�
��7�C��$��-�H�k�!)Q��7���[+���x�t�e ��G7ON�Ռ�9]�� A����X��
sqR�c>�ş��H��˼��^����n�Ijt%�2���{Ad�R!���{�x/���[�E >��q�z��F*e^܎ct���z���2j���م'���cn�%�YJ���A��Mť�H2͊ʹ�>�K,��c-��iP��,���I�8!$�%ߛ>�|��kI����D�֭Oh�홸�?{X5��Du�0�6x�., ܭ��#=�|�g��!s]�"I�K����۠�(�"ME)�Yó���j��_���P����C�<wR�#�T�4�
QJ���
.�S�kW���� &�p�yY�2G���(8�bU*luw�ҳq����[͑�����Z�{��p4,��I�*#Q~c�]0��;;��"��ա5�X����(!ڵto��qg��S<�\!k̙�]7r�:�u�2��ۈOo���Y�JLL�E�1�x�mA��B�v;		L	���ˆ�%}6E�+�oZr6��	+�EI��Dq���Y*�(H��K�(��"���_7�}�����u���N8�6o�/�>�kɞ)r��;�A�H� ��y����|�Y����_h��Y��f����	� ~��'�p��s�׌F�G�X ��M�
�(\���C�d�9��ud��Kڗ�\��2��p�9��a����А��c	-����z�~�L	҈mi���̥իBN�h_$���k;o�/ �?������e�t�A~�<���L7tMC:'��K+��a�b��G��S�\}�k��\��L.�G���ף��k��_�\Wd;|	�z��Px��z�+d. ������i����۲�|�����d�~�)ʇ� >]�&$�x!��~t@e5�G�c)�������w������G��F�M��}(�q�"�ٟ<��8�͘E # �4���i�"b�d�]�NnҠ�>-��8�dp� ����Y]� Hۤ r��	�YX�F��-.go�Ő�3�O���B=ܿ6�jZo�����<�滤Բ�uS�����n�Xs'F����[Y�K�;��kpZj�����톣�P�Vg'���g��FlL'Y��9l���~����w=؇��/	�(=�a}�xҪ�}��R�Z�9�ސ��>21��l�j��&�AE3��� ��m�7���{�n�������xvW�u<�H7�7�
�7����%9?y�������Iur!�<4n���!�,*H�5�܇�Qմ��	���k�$�p�L�Ե؄�]/�>SW�ơ�� �uNO�+D����-�IR	o}0��]�� ��=s�T"�M�wg	�ޣd�@�aZo�W����� �œ�/�s�3������QMÜj�%�i9۶

��1�/⹎�+��_'���H�X��)d�ٰ�����F>��)b����B�]t�2�p�zf�oU3���'�6�����1�q���|��2�K���O��M��wv>�
n;����5a%�ڙ��GW>�8�#�-~�E��}ž�b�8�U��^�qdը�a�no��;��}`���,(��T��'Z�ҭS��g8fV�#�� �ǉv��=۞(�᫳�JK��N6`�m
v�j�8�u����G�G���E ,<��>!}\���~���"/��Jp2́! �j�x�K��	�śq�mZd	�	��+Q��U'}�P5C�Ue����l� |���Ğ�Gi]B�Ӝ��V�*r��=�\�eK�L~J`d��T�C6��@-��lx
j�=A����_�|��x��36��^[� ��|����Q�HP3���h��d�J!�PQj�K*?���Dbn`�Z̊�"2b�s�x�7���0�\��*�m^ϛ��� �\��U�1 �+K�o����x6��`���kaq�Rr�\��$�{
z`��|y�����"3�e��\u�f��2�r^h�iֲk��OΖ8� ?��?*^b=<��t.ڠ8ZP7_�ߎ#׍���A��%�F%v�ٜ�s��[�����T0i4*�E��dKLp���-V]wu��:����؈�3���y����Ԣ\�o�贠�R��EL���B�vI��/��Ϸ�J�HJ3�I�@-����Ҡ�[k��q@y�m��U���u�;+���u���s���J���ץ+z�8����t2���^NyR�*�Ȃ��������1&�\��碕�1�p}R��l���S`���m�H��~�:/u�15ѫo��+^�@�~�2�Z�e�t0��&�!�2]�q_ՠچ��7�lqk�i�x��[���u�ö�A�wi͓�6�d+圩4�(Ms|K����*#�+K:[� 
�gG�4V?%��:ƣ!��U�)z�%����[�����v
(�(O=\;IKT�3�s��X�Ex��w��%�G\�/���icM�u�5)	�I�����(ˉ%|�'v��Y�z4ɤі�e�.���'���#��]0&��8�o�5U1u�Yй�4UH��m~U!�ꖂ�.��"�
�� �g�u	r;v��#����f�t-@�{DA��yGX"%w}�o�5o�P����uD��?+�����+L����?\��L�*�<N&�����T��ǩ�1�@ Q�Ň��X���G}���eu�f�{EeU~�7��6`-�lk�Y�;�����)�uΐ$���e0he�?|]K�&ӡƲ�Ed�|�z�XlwC�PK����r���h�k_�?��巗1\�T����a� ����>,Aw���JZ�Y�9ZKX?�z`�0�����R���@�d�;c<ϽKAZ`��KdչZ�;G�m��غ>�f���R:�ЃK���_,��{*��vm@�6���l�L.Nf��#���Y�H[�XB�S���^Doʔ�f�����C���r�ͻ��ݱP-B��{LRI��/�Y��B�.��T�˔�C����.�o|w����Q��k"W:O۝#�����"C�u�ʻ���t�6�$�X����FO�M���>V�w��^�D}�$B��U�	�a2T��:��@���A�^Il�upF&w��sITX�����HqD6+�����h'��!_ez���>7���>*U`.9 �<�a�R��WH;_�P��5��e�QG}�Sտ�����~���q��I�i��lq20G��*Iϸ�i�rXm�o��*:�>����[rCm�'��y�#�K�=������ �:�8BWE��y��o�$g�E��8xиR��w�ԆI����2�"� P�(��f�p�Cd\OA�DgG����[.%.����i7�
������\T_Oh�z.2�*`\E�E�����r�!Cjo�B��K��b�ѡ�G��cT�C�I�|[�<M�4�<	>F��{��Y������%0U�r��B��3�b>;�7o��`��s��=0��[����@|Nz������?����t>dF5b�.v5�`g6P��ݴ�  [H���L]�cR��ఉ'�B���xň%�Bce�����{��^I����;I�JƸ��}<��:�9�� $�a�5�(;}2`_;�J�'75�S��d{����q�s�i���&�1�e�츫�����fǷw�W�[����X�w˳�!�m$�>k��
NO	���|F���+�*�*k��(���{Y5� �bI����9'�؜X��k\674B@�����#%��V�$IzIivr��E���y�b(<�UK��BHKp������)6���ֳt����»��<��.L�//Yo�4��@} ���P��\��v���{usQ��j�Ҥqu�I�vG��}�W�����D)o��W�L6��(���:����1H|�� 8��O�H.�Ү+�{s��m������Hidn�G57�n��ad���E�2��6�e��ǀ#
VΚ��Jsf����R'ӫu���<E�n�+L[��L�S�i�z�y��$�9���4�I�ײ'ڌ5��S�E1����]�5�p�z�6��"�Yf̦��*'�
tՈ5�'�`ǃ�6� =\Ύڥ��,F N���/-�3�������p	���?
w(���R���������rO"ً5��DW��T T\�-X���_-��KW{N�M���r���~Kf�G"6��ׯ�*R�ȉ���zXκQ_�XX�`�����>e7ַ4�z�12�������Wz�b���<�#��g�Ťy�
X\&iZ��n,dDű}�_a��+���q�G����������P=�ѿE�]!�X �$=fm����	����oK��	[����<�W����O�_�Ajf~��2���mN����B7��祧�2E�W�ŕ>�(����G���If"�+WS9gm�S�UU�u0�Dm�m�i �ʉ�������˺��d�Q2�:W*�Ը���wX����"*�Y7߃D�)ʇ^�*U|�$'�eE�.#���|f�k��B�L���VV��>ʣ$c/qSƣ��$:}�n!�w���&��K����Q �/�ɸw��4}�y�b	E��zG����9l��^rN���C;�k��{���"��/Õ���g����\�E���A%�mHg����J'f�X�L$��skGO<"������u�������o�Q�z�ksU��$A\�wR5	���S1fوP����,U��	���.����@hPذm�e�[Җx7m�D�n��*$(`iwt��/sd��b���J�k*^"!���w�|�1}���MU�q�|���џ�H��}j����hUK>�*�%�X3R^[�T��!�w�����XO;]{�#���+$Y�؟�P��(��[=�B�x^�t�II��'�2/��$4��:r&�A7'`�+��`�����	��Z�s�]��6�ݗ�~�R��o7�އXҌ�n�9� fE�K����<�T��_�7�����sQ~5z�
���yxu�^qֻ�<����"��lt�I�e�;�5ca�����x�%�N��o���+R�\0̡f֪������wz<e���+qj=�%�1hܘ�z��y���I�A*�^e�ⳑ����XD�
���r����&F��h��	��O�8�;}�=�Iߕ��/���8튂������Z��:���3���rG����qT�Y�Ԓ�e�Kk,���&��Q��uzD.�i��R�W���
��k�/�=>_���Ą�f���9��ˡ�c�v)	B���98�L�U�,5tB�a�[�f�D#������"��J ��B�� m�J/��$#Ua� ٙ��,*ƢW�T�~<��}�\"_8���ガ	��  x80��␙%�����[y�p����ᛟb������T8�rIL`�ƛ���@c{0A�%���"���O���@��R]F�z�]S�c>�p�,�,���}�z�!T��0j?��f2���2���	��r0�>J絛���*��Kn�#����a	���a9��_P+'���AX��/"�� ���D��"VtL*UJ?���"'EojD�J���y���1q��լy��7�ܭ׊�氞�:�&pҰԫ��Q���)+��Xą��H˾��ߘ@V	�A���3Nz�3�����˼��ýe|U:\��g�I��ꚤ����.zU�D4�8b
�ߩp~�v��΍��{�k�^y �Od�l�0�7H	K9ڷ��T�+K�*��ߝGT��eUɜ�Wz����)�u��j
�vKG��Úl�ms�7KQv!-*g��/ߝǜ}�Ϭn�����&�H�&��p4��!��	R��U�j�00�,	�kY3��A�-�Q2>/�5D���5���h?6���+�|��d�fF�ƄT�UՔXJ����	�WS���9+�����S
�S�H4��%��O�1���l���1�����|\���R��b ?�`�l�?�]��cI��a�/|A��)�-]O�ۺ/�ʢ�}e��=���҅�>6���M�4Pjyw0�p�ZBڭ|7�����ì/�.��A��ߵ'���,���[�4�,ofH�u$��2�O��B���Z�fM?�%�'�Z?�Ѵ�H&��L��p��H�G��?AMU��JN�S$���'7|��g�,����\����x�d�2b����<z�B�B�6�����!ח�#K��s�a�I�Q���L�vPO����!)�ޖ�z~��V����Uj7�/%��/�)��Jj[ЮɕN�^r I�|k�}(f�%�O�W�d|�w)S�ٱ;NGF��r�������gZr�#)]+�0������U(��=�WU9z#��w�_H�r��9oiQh݁����do�6��L]��lgC����N��DvwS���2K�ތ�ԋ����{��c���@��[�5w=���/%�.�^�8����Z��&���'�N��e�@����۳�(�+��=`L�	���O��B�e�L$��@�� z���E�P��˃�+�D��t1�I��{-6fn0;��ؚ<`�fN�,p��z���˶d�H���PIH�Y�́�Z.nf,.��C��ƨ��yl'{�s|Q"�}_�ir���	�	����\Q��[���[��]���(�^��r��F<����Q�Ҥ�t�#����L��5nL���p&=h��i�J^�ὤ��к��O;� �b����� ���r��x�<z��|O�O�8���wӼ�����o���*ý��X
҆�����j�+V.��D���MQέ��a	/�{�jW�h�����I �t��$�p�G�
�=�,^_+�F@?$c��>�+���R���\l���)�b=Y"��ޞ�S������+،q�*-Ne��~�xU)u"�%i[�<m���
]H��HR�g�9x����mNG�����0�*���ĉ��s�,�M�"43���.
]I=�9���������7	�p�N��,��kMb���K��?�&��I���3�� H���3�b������&87��i�dOC�-��vu���bA���R�)]�I������aJ,���(7C���<�1odQM�esk���c iB��"��B"�j�	���l����Zm���]0��U[5��:������K� )c�6�O�v+3s����)(�puֹ$��Ӌ�#{62��E5�U�R��dXJ����À-
�3��<,v^�1��?X�EE½$�.	� v�T�XX��G��6��j�V������=�0`r��>0�SP�S�������=Ej�����SI(ͨ�U|c"?��zL�o�~�������/Ӊ>��צS�uv�l��-v �qP�d���"��pm�\\>���i^�p�F7=�q�:>������6P�r��&�>���z]t<Il�,��,�s���V����x��ǣ7FJ:����ح����y��ε��1訢z�_����'&]Wc_vg����?���bXӍ,�"v�C��1_HvM�S+��]|{��3��W�Ti�[���i��OP6�hv�"+�,62d_.5����	:�;��:Msn�FȘ%i,��"��w�C�9��un��_�
����,ֻ��T�E�S�ꔦ+�舝��u�ͮ��EͧO��-�9Y��E��o���#-�����S��>�tH��P���n�b� �C�y9��I�[ב#��z}֨Ű�-�3*�o�t@�,�v7~�8ݽ:I4鶸�>=�V�
ZOX�M��=��ݰ5ɗM��k2���^���g}ĉ����k+���S#�py>A]����^6=�'�ٯ'
� +�Gq��	Z<�wq-�r4&.�Ľ���u|ur+�*9r{�Q�T)F�$�"F�[E��*��Ȅ&���{[1�rf��-^�}O~w�����/4�+>������̦��a}+�s`�����^cQr�`t���\�N��H��I�N��3Ã3Fr�c�/ȳ�9[15�q6��RZg�wag���<D�Zzg��-!A�M �~'s��tf��۳3��Y��SL�e���V0���������1�▢�묯��v ��h��܏R7�$[k�z��=��ګ����q�������JP��{y�0	}�6���R���.�c&�?�)����5,z9��Xr��'Uq����>em&�~B��ʰ޿�LCm������ғRJ%�=mJ�A�1H�qQH[V~`y4�y�c.^�I�V�R�Սۥ�-���t ��KC��������X���*V��ǰ���Y;}�W�@MO,�k#>��9�^�g�1PO�3�/"?X-�,^;�:�����f�x�Q�1�Y�j�����c�,��
����/������V�q��ќnN4��<����E�8nM�ߢ��:�zퟫ*X��Cs?���Xx!����k��OWc��3�J��Q�gڀ9w�[H�����Q�zշ����*���?��*�)H�G��ѩ|o�k�y�dEƙ�oCZ)e��^���n�|5N ��a�?�S��������￴��Zi��G�ة�q��tG��-w�I�;�;~��pi-�ej�be?$4���r���Vɱ;�9�����#����P~,Porb��C{S���5E�5��e\BE��	�{��a+!�hp����#xJ���*�֐�Y�fR,��d1Y0��������K��lU>�%?�E�'/;��p��EY�xF]�.�[���ڇ'|B]�§�x�j���25��g')=6HC��&W#�dɂ ԁG��\9�RT-cS.29� ?�Ϋ��m��3w����F*�n�&�ّau��n6����.2�������U�dD����1�hq
�FK僁6�rVհAK
>,��X*��P�k��^GU�hH��_�Z�dk�%_=��Dqu�(t�c�r��d%��Z�o�0�ɿ���z����ΆJg�R��,�4C]&�<0I�2��N��BN�������fS�\c}�]ư>�0�آ�\I�7`D���ߏN��}!əƇy?��v�m���/9�}E=�5:V�U����q7h��eUB���B��8�a��C�ʿj�ԿrXt
+�N�9��ԂE3��*�
���	t����k���ǋ���X�J� �?�Z*�l���#:�h����!~��k<1��QB���>L�DRB��Vh^_Q�&�]F���?Q,.���\�&P ��G���u�,�8���)@�q��\W�ft�s%�ui^.�F�	�un�y���0�1�p�[���Ē�����Ѝ��4��VhJ��5��oT,W��-
.���ԥ���Y�߰sXR'��<������T �I�0:�z�Q
�O1�����I�n�+�`�+�:7�%ٱ-7�Q`ik{n��| ���8=,I��:�nu
����M��7٨�L�C�V��M�1!u��7�XUr��H��Ϻ��6�{荌�lQI�k��{����i�!����E
���}��F]��?4{|�E�@s缼��4�XP���W'T�BP�3�E�U�=aL���BY��\r�p��R��&��j�u�22�~���Ϥ�P�T d{K��{Y2�~g ��%o�@������O��,?��je���mah�ԏ��W�g����,����i�T�ws:�����|����c��vb��	)�)��W��׭ɶmZ_��f����d����C��qL%��d��*_�Q�b���B���;��֪�q�p�A�MSn�]��a��S��&�����Nk1u
���d1�g���ثp�:�����8��W�Y�}�d$ lmպ[�ga�y�Gs�[M� ��8��.�ڝâ���&R�W�A���^�rFJ�3kC���!�Z����QDJ���#/�@)�6;�|I�
ԋ�����p�ϟ��B��\{[��~Fَe����&;����?v��1���(��/��Rc���:8����b��sa��o}3�ɔ�Ժ'����1N;d����/��+���7$�V�ʍ�{,�����`jД������Ǫ��B<2
A�y���Ŭ[��4;^�ux�CŔ�Z~�gq(���AL�KyӁW`�G�N�gֵ�@T,Y;������|����#\�&鴠�*Y���������,��N#2vNx��j6N�%�&�����m7�6���1D a <��ڡ$���I���q��S�6f�eE����%��1&WVi �9څ��XSL��ιnϋ��А�A� ]�����T���PN@�WVj�%C}�g��?�!��[�@-�T(���y�lan�!CtO	��
M�X�I�]�	��4�m��u� �n�%�Q9��6����o����Dw���x�a�J"CE��b���6�v������
�_ݨilz�	�5��n� .�Q��}�W�j(��|��?L�5���f���*8�@\ъt�O!���9YJ,��ߍ�Ȣ�v�8e�� +�ߴ�K��[�R��r��]��{>���3�h���
�T��y%]s�P>��-�>�;�k�d��4(I�TB)V2Q������U 奜v�є�lbȺiK<�$-�V��2>����&ac�H1%�a��X���\Bk$} |JUa��y���
jL?w���+���la���h�c��'1C@as�}�3	|+i�
Q�9֚�ض�
)�ޢ1[X�ٓ�:efb$4d@�.��d[��Lj��.f	�{ ��-�U���(�I/ɪ���{�F�/�3���.��odf,?����I���c�+�;��f����9�yd7{����T�W�g�--4I*�urb
�ӘKO�n���!Y���x0u=�J�+��Q�^G�%���!/��D�O�u�#j]��`9R�ߥ[��O�]@(�[0�i�.fͼ� �w��57��K�VP�4��@���a�ai��y�ÒM��f�޸Q(<��㥯��ӑ�����K���긋��!{Q�W�Jژ��1k<�f�)��.�w�Q�
���v���myw�O���lح�w�u��;m&�Ad�,>*���B���V���R��[�$В����Z�������e�ϐ[p<M�~[����i�~q��>اxZ��愃=���j�m\�(nڧA�,�$=B��j�?�C���;I@���;!�S�D� ��H��.�Д�Y�~��@�� >i~a�2�T�]Dai�S�z��B��e���B�?g%	����J$ލkkY_�7���+� ����^=��
�ް𷯛�)�=r2w��v��qŢ-���CD/ȭ:3��ʹ�m�Xi��ÖQ�m|x�L��{I�a�u��8�&�B��bPPD�ۼdTyE<=4n��X������q�[�}f���?�R�_W�h��/��)$ℂ��*�d	Kp�R7�u��lC����.�������@88ب�{��������|p�(,]��S�۶ձ��Q�@T$��]��&��ِ2��l3h���0D������EED���׎�!�dy7�y=7W����mRR;>x������-�r1����&��3����i����b��93r�Qq�yح�h�)�uKj��7z�_7�,�H�^���6��ؕ�k��N��LjL8�ٶ�G�4�y��?&D�WÑ�4v	�%+O���s��I4�͔|��64�z3�Ѻ�s�Q�jkw���u�,���`,�(2�����I-a�F��P�2��k��s#m�H��;��z~�ۣ��=<��XT�WE�4�R���P�Ow�׊�{E(��{]r�Rg�:���qتR�&z��,�}�	P��	(9Hi�Yc_^�h��w��ȵ���j��m����^��l�'�i�S���V�1�!H�R�P�*O���\�m�J_��}��]W!�^�����!��cI]|!�*���>':ɷϫ�!�/�"����n�º��A��0#�"�S �Ⱦ�7��Kh:�[����a�j�Cc�|s� ��q�pR���0�\�A�ѭb5�����<��U#�wR�X~�-�Ӛj��ε9����ʵ]u|��%��@���'$�E�栮�����;8
�����h�߫4{u����0a[K�E����~���e����ǹ�u|�p_�m߭���Y��`�/�w�Bu,EB�v��x��M�z�wc�ǓZ�7��n�M9(�7�J �v�|��	��=��pks#��J�a!��U�y$\G�,�;Hβ}U�s���/��=��h\V��V"K;��L�)3c=tzڟ)C�ɱ�����n-P����uҲ���מz��z3kk��I$"���#��#5��p�W��}�5㙥"�UV?��>n3i���^wf�
�QC��1}��]ق�x'�����ϔ��ߐySr�=I�a� ���*k}-���Ѻ!���NB�'M�Ԗ��lk��B�I�6�o����qs��xS�g�E7�R�y��mˋ�����?���#d��`�y��҂"�j�:�Hm�*! �m��1i�����8fya�ִvX=^ϋ4��|.��VKMoS�0���*}z�"��3��e���X#�5�j�@*���l-U�1i}�P��|Q梧O`��&��bY��ޭ����C1�*�@��xȖ����dcW�f<P�1ҩ���d�-�?N�n�[6 Mh*s��m�'S��Cˋ���LIY��G�~�@Wb�����gj)�04J����:Y��)����=j���?����WV&7���U�$A�Av�c�e���F�T�O�q]D[��'Z\����6�����R���z*��a.k	�yS+D��#Oň���x>òj�B�yfؾ2|	TY�xϊ��2.Ӆ��.�Ӯ�=s�	���x�R�����o���|�C����wu<e����yg�nM�6�1XV�g=��|1�
o�=��<8tT�n 'R��4��e�Ag��l�w�G��9�;a5%(�x�F���aہʬ� ��i�:���,�P���L�m_�j�TV���A���Z�U4�Կ�e$��ԋ�:��U���"j���Έ5Rn�b]9�#2x���
s��/z0L��m�~�M�7E2!f�zA�t���f��cCݵ�|Ce���� �G���a��.�pΤfz	�%i��$��	�$~�e�����r�H=��'�ΏK-b�y�����V�t���@�@����;d&�J��50D)�ěJT����#��z��vp�3S̰���yk0���)��b��D�l)�� n�_�k�������d����v�(V�i�IAA�0^a��op}�>
��E��|�l��$%��ӊs6�������Q������-�칾��Y�2�Zd�8�_XРtm�Ԡ).;t���=�B���=�����`ث�~m�|�����uE��ݓ���ۀ*%�mU����
m��}lPo��L�(�}X�����"bR�bS��GU���\�U��I�uW���Z�>R��pkl�����w�tAc,�o��0�x�W9��k�Od��}��|�2�k6���v�&P����� �&��[��g�!���
��E�"���N���[�{��l�ˋq��ku}�|CrP?�}���:�ף����v�GH������ig�5.����?�� }Ӭ�;)}��/�W1S��S����M��O�\��\�)O`�+�vU_�|�_��>g��F_$Ώ�����VQ��y��^v*�)y�k.��M˒�󳄜.
�r/ю��ח_���4�����2�w&����u��Qkb��Lb_���|ˍ��qaN���~8-GkIv��e����O����\��]��cEJrU=�a��f�&dC�&��>^[^7�pXvcf1�P��� �Q�Ϭ�&Qố���Ď�@+�Sm��/	�F���Oȷ�[¢��>O�X�����l�\i����01*��3T���&�:2���C��Rs�Q�� os^Vt)k�jõ�N�aAb�f�ƪ���kl���>�Ӓ8�/��������t,��E�l�RN�)%N�z�"X�?ng��,����,1�(�Z_o"�Zz�E��;��~	�|���O�4��� ��T�s�	9����)�l�	�j�# �^P>'a]<�%���7HR��S
f�� ͽJh�C�?��O}v6���ww�Z�g3���w�I!Q�1����BZ��*����E��v�M��+h?�A�U<C������ҟ��r����
�7��'�?=p���(�ʥy$kQOk��yc��냿X8����(�L�/b��	ƾWk��?�O`rqO��k��4dn���x��ِ��2ᨕ�D<�4Nf�.��+���Q�TC�^;B���?��h�0��p�iy].ɔt`�5㤙^�)*]�k��C��L[e~йy�Pi*��*F� �2"8]�S�;*7�]��"���/M�-���?�,�h�V	�`����
�O�{� �7��T��uȮxy�i��t��J�h�R,��&cI���&�� W6w0��x���>m�kv�_�I�� �Յ9��3��Iɷ©W��#׃)�S�9V\%R�ZЄݐ2%O�\�P�![ME�n��AY�*\��Du�����O /#5Äo^��z��xЊ�7�=�����;J_��ZAso���z� �N�,�v���w:����r�C���s]�uR����8�۬}l#_xr-98����a�UB*��y
m�'9�a(��]�k�Ӑ�
��~���_��r��C%�ӗ�Ye0m۾^�r�o���=?�;.(�,58D��*7n�0��{[�������îru�`������r���%�f��ę��-�
�b�'NKNUU�
�������MɌ~J�٧CY��1���M�y<��� ?0Ņ���[f�0�up���8߳������6��F���)�?��'��r�T�f�WD�]�vI|���NE����.n�I�u�P$�i�T�3���a;�h�l4�6�!(�N���^�F���v�*�<�ɚ�3m=������y��k	�T������l)P��QE�*s�h��b�B�l�k��p��V�Q�L��h(�����01C���ʒ�ԇC��[Z����Z���y�$��&�jF	X�:�=���@�<��W��@g��F�A�a���s�1*��ק�n��&�����9kj�	���d�� &g��p���=m%��x�}?�L)�	�ɲR�I����R����&%j͟I��_���@���WV!P�F�j�9��D�B�֏�<ɘ��o�K� �]�5�
��fCn��ҩ�.7F�r�L���J=��(�򑖗~@Z��q����^n8�pH|��Út�u8�Z�^x[����)ٗ���?]H72R�|R6���ݐ�t�����%>%�E#�YV� ySa�	Ԕ��.�,y����(s�
��"���jͲ�Cc�4�/�m�~d�IAV#�����&��VWDɝ�,)�2��Xkt���TE��DXT��G,šA`H����G2����|f1#i�)1�e�W�g|�tx�����f.r�Q$����o�t޽%�n(������~�n�9{s�/j�_�h���90�����O6.�#��Vۍ�,�����4��&%at���l���G�R��y�{�ኻ;ݔOb��`h��RXqڢ�S䖆?؆���)����sC�4��%��5�7$6&ޘ�L_��b6ƕ��#^�BQ�9����uTX�%� 0���c�ng��l�"O�W�u�e*�8 ���s�g�˻�G����Y_9���"�0C?�Te����_^nx�h9��O�o�kw�"w�E����q�5k��݂y�O�y%lť��֒�v�+C�/5�C�$z^�D:*���{!Xv.�D:�����82�.�T��o����8�-_R��7�l3��z���, 
�Y1����|G��8*�iP�P⩂��!���n�#p��}�+�]no��++��seu4�\���S����So��us���&i^�V_?�����1���]��e٘͗�+;��M�vH+���aE� �NRJ�Q��m`T!��`��n�c4�3*���8�����.��:�\�&� g������r�Ȓ7�'6���r���w�R�G���o�e�/���?L}�?�K&O�yt��B�~CȇAu�:�\���>Sb}3T�m�<��A=�&Рv���n5F��E[x�D]��:+��ϝ����e�4��1����	˜H��5o`|��
��ͱ��Y�[b�rzG0�8�4Ӊp+Itj50u��jv�|6�A�<݄�*�YH�u]|@,Z��E�T���� �o�s&�{@�U2�/�RQe�BƝv�u^���:`x ��L,;=��>)ϵ1�h��0Ņg��O�-2��+|�����QZ��SN�o�x��*��Q7�`���N0�5�������Q{PD����`$������zV�y���V�՜���Aq�J|�Q�Oj��L��̌���������_��(TθQ�F�Ŧ�Qv��GkA��	c������C��N��DO(�V��/�0Y�2<����o�$��Y���oƩHJ1�hb�}�N}&F	D	�����M���n�Y�Bmx^�쩬�:�k���1c��4��#�w^��Q#t}��j�Kz��HQ.��`i�ϵ� �E��B�"�+]��#�`�
t�������Y.�������~�O^G�7��߆!t�8���T�!�N$@}�Aԙ���Wٞ{���*�'�DsT����6��#p������|�ID�
�j�8&&�̚�tl>+�@�\������{2�Ĉ��f�	�=dU� _z�6������V�\J1�m�w����L��&��Ɔ�ux^QȤ�q�Sz2��Q��� =�z3f�u/8	I�37y�������
��+<�"��F=�r�|��3������t�'�KD����P��nKV�N���s���&n	��"�_�;+�f����ӫv�i3V�8�A��둕�z[v��ILb�nѕbY} J�XA8�"����^����(I7M�x�̕L�X����O
�7���a���K�-6s�_�Pa�bAj����++����.^yK�\.�mx��[n�\g�R�*�O����w�ƱCw� .F��fo4F�c����-{�<��[�F.�&�~��po]@1��S򧦋X lJ��P�+d�)	7���#D��/	W����
+-��N 'Y@Z�B�u�k%|�)�w��v��.���Un~o�����Pn��K)L6���d�	u���v��G�s=���8��/�վ#��#�7�s���E�ݖ��}� ]�45�ã��o��X�NQ��x���k"Ws^�����c�q��z��Y��m$Q�����0h�	̳Q6cAq�� $���p���B�Xx;�??�fsuq\�\lD�B������7��(�M��U�@���GՎ��f��=t�.ḽ/��f �o�]_S�Q�̉^I+���@�H:,��	�Wڞ`�5�P�gM�/�%O�[�4	/o�rc�d���:`�-\�2�p�}6}��Po�qI��)�b,&G~Lm�K�W��~�����v!�jjmx�M^�\�1ք�Gh䤐o�^�sV���rX��b�����A���'��\�P���2�����6���`����#��W��#�,$M�f���/�?��Q�;�)�A���怢a���h:����TC�8��B6�R/�Քc�s[��@�Y�x߰A}���\�U��ڗ��mq�aY��������o�/��\�X�R��f�y�HS��}1��ܩ�lקoP���h�7�o�o���j��ǻ��	u�-r�oSԓ�k),��W���WI[�Y�\G�?��C�d�^fX�8D��=+�㱹��A�7҈�~6�)�'�t�X�?��A�O w�Bᐿ��3b���e�Y���_A���({Y�X�������L�+~S���4��~U.R���Y�A��:���S�&�^ҹ[�$�rj��黝���p���~�TT��;��#�Q��S&�G�<����<�HT���f����^^��>��SuH�!��� )�3\��9�3�A�F}t��q]{l�̥F�������0���QH�59'#א2��x$lw�����s"���,�Ká�>p���⇌����r=x�B;����7{�Pl�4�\�����j����A��3*�l�-�f��� �w[ؕF�ѬPB��1�۹`��:D�^�ٶ���f_���0#E�?���Dm��<�3���=<HW�u��9�iu�gj�����l���<��Aa;0�.^�
X/��q�>�����}��l�i�"�����$M�]�|93�{���L���-�1�[B����#�zz�ぢRg��UU�I��%X��5eDK)δ��Rz��7$�E����6�5��g��;���~A�ˣϡ<�h�n̕/K�GY�	C�i	-MH͉M>gRb��zWjU���doR���';�K0���#�t��BK@�<.+1&>nb��-�N�f����\���0M
=o��f�*��vO��pa���mHXq���Yw�j�D��ѭ���m��&-B�]�^��8�Fy���Cn���{X��::���x�/hqC����dq�<���`�ɡ��yf�{\��黯*(�^�}���Սd}o5�|e0g�Z�=�����?�����������ñ^�5pg�����[���64����F�2���c��9�l��q�rc��7�XbBm�"� '�W�4.��g����̎Ա����jC4s.1罊'��8�Ǝ���4p��*�gl��'�Õ���k����-V�Pﱔ�DT��Bg3��h�E�s=���u�M>�}�*�£4
<.r���W�g:<������UF+9{�D;�i��zq��W ��+qC��bk1�'7�9���;TQ�v�d�4�9
"����K1�O�Y
`����W0�^(Ջ�M���(��^��� wdvhq7�?�0r��}�'�������<�xeEGE����6?��s<�W���WEQW�BP\10+q����达���^~%�sp��Y��a3_����%lX�g�@ �ԕʖ7��t��{��P;آ_u�4�%Й*rd) Ά����l!�'ῳ���ꨉU�B{�Pq��^�Vqb�qz�\�U�`�ۄ,�w��1/n�-�q��0�D��!q�H��)�o�6�o�����Y�A���c�{�Ǉ�%&�&��獄�A.��`-���O��柳�����~lG��I��z�n����H	>�?����$F
��,�n�4"P
�SMF����3��L��]���G��&̊�������P�Fv�]�6O�����AWݕ띬Aq�\<q�� ?�S�=�=�+��S&�*M���#�5K�����zvݲ�D���f���V�������y�eٲ�	�%o	���y{�����⁜0O�9@N�<S,˴��m�L؀�p�l��pq��i
�?���r!�w���|��E�369;�͇��<�$@� q�8{V�b�_jt(CH^`��'�A��sF0)��px�o��sA�H$�!�TR�*v*i�i{���:�����1tO�}r�$-"�0��������=~u�OU(��2��>�0-��iQ��x��Tc����G>��D�z�`	^DO�X۾J����ru��T����a0+I��l�T�W���-$��N ���� �r�n�j�D4zn����ѫ���c���Y����k����0��5�����������vϔ(�{Y@RY���0����oS���|^�(ĸ�4x�:t0w��
�.��*���٨���[#�����_�����?��7�p
&�e�a�Er#t�����^,̣{(UH~����,���F��A�9C"r��#IG����j:���b��?6C��e(hi�P��#N�������!�~b���t�'Uo]���vc{F���t�6����چ>�?��|��fv��_�n'��.��~�
_��T�zq��Ι%_MRܼ8��0�Қ�	9�Gt�~V��%+���J�4צ3�TҎ�Y�)�GW(��[��I�֮7k�bTGϙ'OU��@���ou ��{�M����Uu�Aj?�/����D�5��7��T�����͠�)Wo��$�8`��6�7��פy�f���A��TS���d����I`��nj^h�+�l��}�*?Ê�����7Cu9�B�o�¡��β�}�	*<n$Q���O��͚��+ex�alW��V����sv��t�o'��
��wy��ă]{OBg���L�ڛ2F#��Gq�sϜAu���T����R<I4x"�::_�g�rc�ʤ#�%�q%Z~<����#��n��ra��|�1��2_�����7���8ZJ@(G�E�zk���I��sUT߅���^-�,?�ݺ�4����B��
�����[_�$�&�ߒ����"��"g�W���;�n"�U�����rGM�aA�%�A��N�]��+��N�t�ύ��&��i,?T{��XҖ��K\c�Յ��ɖlr��D+�+�y`:2�xѻG�\Zu��B�z��{?�����$9��}��;�|Hh�� KT�1�pC�Y���PN�ꏆ�T7^�������ܝ8+)��9'��؊�t�
	}W�9e�j�[nF�'(g
7D��?����om&�66]~�?B{(� �x�$����*�h��P$J4u�+߃ݏ���K1[�v�8��YL<��gO	��	yK<\�#�>�%hV��.�lG��S`?�OW�0�l�+U*��ɽ��rn��{�)
�q�桟�6���@���w~�}�6��r�3O�6F�)cc���l�. �e���MA�^�T�+٤4�s��:��R��j2�
` ��ुP�N��4���Sy���E_FR����[�I[Ѹ�<N���8)�d"��sݺ�k�2
*�b��H�T���iԂ�L���ռgs�ts������w�K4+<+������9F�X�_�3X���0�x�zm1bd��&���R���v>��1J,���z��x\t�ͷ�x�
�����RZh�Ye��k���U�%,�oh�T�s����(�՚�*G���-��ʨ�4�ҊFt���q��F3i�9)I
N6��:dL���U��$��<^|eV�^�>�h| @_y���D����_���P5R��'�d�k-S&�C#�X�m�3�p��[D��o6����CV#�\�J��Z�΄%��=;a�Ӿ��6a�Py�
 �Ӵ��zZy`��:,�Q{�֕s��jC�;�ƴ�C͋����Y��s�G��.슇�����8�8�\�lfs�����޶鰄?����ğ�;��	�����dP��l#�����gXg��i��$5�j�-��:�t)H��m��7�)C��"����D��k��%v��"+�iUծ�ad������=��*L �K�˷��f��O��ؤ<4�˙�kH�7���ل'%��a$خ-�g�y�E*�QY�-�����9���Eғ#:?o��3��Ishǋ��l�%�/Vq�2�O50��6j�ލd���uK�ཟ���Ao��~^�7��-��hML�����>$�%�Z��g�V�|��~�2t��*���hA�:�5�s���pr���I�!��q�D���K��0>���˞� �g]J�����z�Ԃԑ_� ��ȧ]^fNw����y XYό����vR��^����:-�!}2`�H�M���qy�tk;z�z�R�a���T����1�P��8:��s<h��a�yr&V��	8X�.s��`�p;8Q!Q��|/+�0ޚ&/f���ZY���#�(�@k@h����pГ�ތ~2���	����&��8^tN�<D��:�H>g�V��D�ai�@�l�:��}]ۉr�2��E���f��CF�����d=�e���߸����`�8ߩDqԽ��l��V�\��dt�̣�hۍ޿`�A�\����+�	ٮhk���o�&�B�2�bd��h�k��?'��sX2��.ԇ��H
r�<zq��d�q����CWI�"JE��+��iP�r�I9�.I�\�J9U�a����>T�2�n}�a8��W�J��x܌��l��e
�lR[qGO��q��>T��a����ku�� 5���ܻs��#�-A֚�
uv4�a���Ax�nd���pX��nt�,���UOM�)�2��>}�z"�tH� �������QZ?����S�k�T���c����.�!B�J���K��44�$���g��+����dQ/�x��5ybWW��!\� �揳��ד�Uc��уLfЪ��n����8h��Is$��t�t�Cwǝ��K�Â#fc�f�w��B��cZ_,T�ŗ���3ͤm��_�i�Ī�T��,���~�7�fw�b�o��&8"Z�>��+�~�����&(��A�H��AO�hpEB'��ϴ�����<Abo��)���9{�����8g^�_�����0�/ڏc}	t8�L�����j�3��C�g�\nĶ��0�Rz":y�A�U�
�CBĹCG�W)5�=�X��x�_ƞ�x�u!�Rs�WĤP��3=_n�l<�'am"���?�#6�\�q2N_�r� gj
�.�.�ݓ��x#�F�x
����hh}�E5��/���]��������cf� �B��/����1�i/ހ�3���&p
�����,��}.�I�|�A'���[�-�� `x^���
J�����#�)���]����(�F~���7:�c\��"�~Y�d`��~���%���kU�x$rc�n��9������*�)oFm����cr��a�9X%XnR�}�2��~?����ҭ�-#V.f�K�̚�����=���&�+��з��.��=�O鲘�r�����{�Z#��������ߠ����3�trU/���yL���6��̈�&bn�~8���Z��N�T��)��
�'y��V�c�+��{�����c�Żٽ��/Ɨ�g�W���(��T�~1deXc�
����w�?�Fo�/*`����(��V]�;s޹e�H����Ө��tZ�g�4�F@�F����|k�'������ءI�K����M]�d��;�Ǌ��d�>g����̕B�D�m&)�XU��l2�:�������lEBB�߱�6�d�{�k�[:�h������j( ��AH�  JrC�/ȫ�v
Z�q.�w�h̊���0(C<��U���SS���N��FE�E5ȆΓZ޾Dʚ��H�&oY�SAʤ�Y�x�.��?��%U�t~��}U����r��O+�u����:�A�$�B��2�NR�/�,��O�kh�Ǟ������k�椇��!�V%���HpU��D��V�N�Fd͎�����H�մ��_�څ����3�0��+�?FT�m�M��$�>�����~ok�S�=p'�(�����K^<X.+����]�o0�s��T��t�Y��o6n�,a����E�K�"ϴ%gU�}���C��eB�e�Hb��M�O� 
]^ZnS�B`+��M�}��)��n8U8H���%���1P�-'n�]+;�}�a�
H�����uڗ��T1�����{�]z���	0~8Τ�A8�p΍x (X�ߕX�,/�2���Is��*�_�����"2�\w�>ۆ��	����hR�U�V��=�ݦ:+[s��^,U�sH0Q�&���@M�O5	&C��D�1�;Av��=��h��W�Hb�*5�
�d1�U��a�������w����U�e����^��!D�u���u%�W�K�O|�S+(q�&c��iLiDL���3g�,��6@�:2���Bb�^4�O��[�z(J $�gQ�t�8	��<US���e�'�r��Y�s�8++�
�A�" �su˿��>(��Î�1/E��߯���JF�?�陼J�ˑ�:M�7�5���O��!����ɰ���P�5z/ք)���z��)�L&n���s�"�+��I��Ty�f��c�-�������	+��-����{iQ\�ݜkY*c��l)Ц9����ԝx�xu��>�ӾE�Mu�膽�0����Vi���ij>X��j����,%��dUkW��|�۱����=������82li���XM:���'��1j�'�ռ�F*��*;W'B�d�K��D��O������ǰP6�5��0Q�
�����C���,��wy3�C#���)�J�����ع��(�R�,�Ӂ�;x������i����v�-�M�tUJt>�#��/F���!�`�����_���0��	�g�E�'��DC�FjK𙼩��~�q�N����N~K����m���M�I>>�RQ������<��Æq0�Ä��,��:`T�wD���>�J���DS�\MQE	����ځR����~��������:υ_��W����]kM�N�+���d��BM9TYf�癑:�w*ΉS��I��-�IyFkL�c�i �s_ڵ�Ķi��NE���A�X@�$l ��H{M�U�͢�X'�z9����b�o�)/��7�� �9�����:]/8��P���FkWKv~�Ξ�F���*��ihn�l[��ew4]����@}D��#|��V,.�3�(�d,hw;_0�M��6ʹ�����@�$��|(u�M�=�:V��H~П��-ؽ`�xJ@� V�ʣ��[+0[Z���ʑRu�#G<�=Ɛ�.����3m,%��4O��i1`��G=~��\�%^��+|��l�&��������Ի;J��%:���A��,����{�&��-D��X0˻���j�Y���2  *Dx-5�x�B"��IB6t����賏��s�4�m����ͪ�~� Q*PBn�1�<��3��1�f+Z�m�_>�b&7ޥ�����B��u�K���S_�c�[ �~\j�S�Y�{8 \]f) �����Iȣʳ��l���	[��#d̢P�T�s��� �l�}��H����l�epJ��\�y&�rkZ�m*��<x}�=��s�|ge����Kf�k���Y5ګΡ	��	�6M|�Q��:�}���t<�2��(p_�m�d�����n�[�g>��fH����__� ]���Ɓ�;�f��2X�ꦵy�Ԡ�2�*b�a3�����l�8��K��s�Gbr�=�@(o��E�b�(����RW"�`x�f��7�\0n��Rs�F�0�UȺ"��cܐ�%�ݺdU`>y�1"�"#��>�i�1;����.*_n)������� �Iu����[�����JqJ��`331�Y��3�a��~)�D��߶6�Ǐ @��7a/Z�1/O�8�mEe����W5ؑ~/�8�ϕ]N�'��K�ϰѬU+�yV5�5)DY�;0&M�7�B���A*Nx*�K��y���IA�mb��1~����[��25	��t�%�h��`;~����k�����Δ�9	�fZ6rI]�ޔd��2s���eզ�|���*/��TlLc�)�n�&2;/cT�7���FB������T
gh�ҝ^vOQ��B�;=��*-���G�$��ׁ��/{�!��YT�ߍ���?Fɞ)�Jg�/<[�v��+.��I��NG�,հY9�1?/��Q��=X_��k�1礗kT�[�d�JȂ��2\����G�k���Y\q��1����4b>�]R���Iޡ6�
^�Z�<����3�pK�!z��>à�ʞϛ�ҵf�J7��e��ҫ�H�u^;Q��d����+�o��Φ�p,���#�s��˫Z��_ث�1:q��%�>��D9h]-b�~qѹ�尤�fZD���I�o�mZ)x��e�\faT�M�j���J$b8�Q���,��D�z�c��G3��M�V/�3Z��5^��'>��=�1����C�S,��[�qi&��*��v�g�8|���:Tn�F����*Iy �8���~T˞���d
*,��b
�l�FŠԍ��JC�U�p�4ا!%nʳRׂ����X�ylÉ��Y�����K�]���RN�b&��?|��rC�̌����_V��8�$��*|ް�}ř0w��@�4��d��,��5ޑ�r=�Kgi��_��.𩘜K����mٝ��8�[Gg�,c^��ֻ�P)�K�*ˎ���Q��>��U4?=ؼ.@hk	�;�� yv.���wD����R��)�L;�X�p���=�{���<���F��uS|w���ї��C>��"̓&�p�T�J���1I� �{C9w�h���	-������%Z��d��f���!,�%^�>Ե��� ��0��L)���2���t* F6�7[f�3����/�'�LB�T3��&�	Z�e�+(\\~�
�[�n�*.����"|��F>�eg��"�_��Ñ�"��7��,-h��ʓlj8��J
p��+��[(�X=?C]�GJ$��:��|��X�uIfwv1����t8o�l^S�F0qr �6>��dO�
����UՁ�*p���g`��ӂ�����/�u����m͍s3�#�M�+��&��ؤ=��I�@�o�.uk8���@�� �uK|��\��M��E���%�Y��Z�k��@�<�\���M�|Z)!2��]��C$�*֔лAЭZ9�X=�_q^���>��Bj%�`?`�r��nՅ�=�b=�P��9�M�E;����\��h�?QF��z�l�;dL��rid��$�|z�6wʚ�� 8��GQW��;"�R2nW7����hV�a4������{�iѤ+8R1�����d�L\������O��"�0*R�pt���gfՄ���*�
nx���������W8����nv�#4xEf�L�K�t�� ���UI��ߺ�o� ���H䰘 V�%K�;�+W
�z���>�����<z�&Gt�:ָ�q�=�������ь�Lg���/B��P-T�����~��?}���Tu_0�J!ۧ:��~�]��g?�.&�F�A&�]��m �O�����[�O�4\��/gC|�p���e9j$�ս�(��Ňr��>����,���<X���	��RI]�=m�	�<�ӨA4W���d��2G˥�-��Z"(�BH��%���'SmbY�z��4i�R6'��tK(���jt�?B��N%h=OQ�Q
�?f�#�+z#6�f�&�Y��B{,.� �b��\���D�r[Cb�UU/�� ���ut1�K��&bt6ޱ�f��G����&�m��K\T���G^U�����خ#��;D�C~��6������x�Xs�l�6�ģ�6�fb�3`�Q�<�3ˀ4�Q~���/�F�B%D�#6m�2zv��gL�S#9����8�P�e��L��3���X�oK��̢Y)s!�|"xU���?0�����Z�; ��l�y�ҍ���L ��-��V��_�CL��_P����l����C�n'1>5^�{�g)��	o,�Z�SV�����W?���X �����p��I��������*�����6��X�%g�Kv���<���K�;AO�>� �8�/�����U�~3���ǿ e��iԑ��f��j�������Y9���Y������K���>?����(��]&I�g 
j�7�a"���p0_)Wp���"�LQe�fv�ð/�����kD�̇?�v�A�o��	�=}�ӎ�9��Z+�����T�E��K�~
�����c�Y��莛��&\9��lr�O`��w�SEj�@e��`�ް"ԚH��{�;�3����rϔ�F��jA���Kō���@/�TE�u+@��픐�a�6�\?P`�OU0M����N�'m:W@7enїy�j�T��2�M��#�5Iu�_������nr[:�w���`��A��իX/o��r
�����'bR)}��YT��<9�m�nB�(�bCm�_��R�?��;S�s��C�!���%�6-�"lTP3-vM��q-�S�h9���>����@k9񱧐B���:)R�g��u��A]괡�U�fG�F5���;����\=�@}�{����X2��J�$?O����k���UHw�t�
����Y�E�޷�W�?����y
������[C��frP_&	�̠V��%Jl�:^��_G�v�z��	�ަ{�=D��'U���/�F|��@o���mA"�jѩod'���4��
�\P|�`�*BQ(9��/yln�w�����UĹ�?��'�B���QBL�.��}�W	���Y9�a��yhB��w�k�`��� {^چ�E�5.=�G?p���wU~B�/*� J������W��'"9M ����$��1�cPv�� �$��(����~���� ��Lz��-�=˼��F	�0n����W`�w��v�+�+�~(�_1��.c����*�饩���	�sAݫ ��dxÈ�`H޼�&���S�Ex�Q��^YF�g�KΒ���ε��z�A	��~E�sfo�HHaá�'
`���9��#��` m��\j�}y][��d�š�le�|��]�q��"I�4X�'�\O�P�-B��"<7⌶�D�����-�V�z܅.����m��:O	P���9�Ax_���^��njz��2��[�Qs}������<}�,W�����0
4�j}lB�˓Fn�Ǥ�:�T�.���x<��9Օ�|�i�)l1a1�X:�X	p]:]�f�#��nyvW�ʉ`B�Q1��h��t��Qn��t[ �j����b�N�>��Bx(큋U�i1~Cu�����H���9�hn�y��,��A2�˲l�BBUg����1x�ۤ2BC�hcGKqbR��0�z�Y$6!�
ޠß���Re@υ�?}��M�ǂ�+y�\�mJ�����3��Zk`����Y�V�&a2�����Uͅ��d�D�(�Ps�/Hy�>��~�8����"�EΜ����̻�Q3��+Rݏ����|F��o���z�>5�$G��q��(�>����M�"�kz��	����,�Zuի��
�TS��h( e&"Q�Ց�Me[2u��>�� V_cQ^}�'6���4��_��+sy/vp
Z˲И9t���4F�� ��H�{���j����ƞO�C�P1p�/T&�yzގ�4b�C����mΏ��آ�4D�h&�g:����Τ��j�bD�Kt�����ξ�DOO&S]��$�p4�5�����Ģk���X|�C�Y�&X�b��V�73g��t7�
'�M��ߺ�=��@$�h�oW2��ٚU}�̬��S[iZ�>�:j�qwh-}�^�}�����Wg$^3�(���j+�h.���F�d[u�ҧ�~4�B.����J1��H'� �ORʕ���{@�Lԕ����q��dλEc_�6M}��1��@b���P���gD˪�SBҺyVO���u�>�쫚���/:�T�w�x�Ԙ��2��R<��5a(���%�G���^!n�0�"�jY����;S)�hD��W�f1�fx�fA*��J�j%qAC(�% �X��o��� ��M�=8-e^�h�K�'4J]	Lֽ��e�[ʵЬal�l��n@5p}���T�D�� �VK˜�Ҿ�E���������jE���+hJ�)����O�)�Λ��
<�E����\�i)E��Aػ�Hc�᛻�h<�zx*ӮZPV�zp������_l���VZN�u:�8�*���e*��r�Z�9�����Ɇ�����[țm�&#���A�S��
-��*�Fȥ,���+u���AE$�t{���נ0���p;g�+].3�@�b��y/�wy4�f�V���j�M7C_��Xrs.�z7s;���%�D����)
���\9t�*���+����Fb���j�JP�9-��Ū��+���_T!�[|׬��B���*�G�)5f�X��a%iS3���
��!B�v%m�CzR^ȷZ�T+X��D���*2,�eA���V9�b!�IS��a�XY�9A] "��F<�����'�ި�P)�r�E�"t��P%8��^d)�!��[�{��i�dX�?��wZ!}k�$`��N�4V凣;�Yy��s�ҹ琡j���������)bK�T�H�t�C������AN誣O7-�O�D��������;Ji�����u#�[2�f[K��>�͑W1VZ��N�������@SȇO2�����C�1L�μ�v�]�>���V�A��b:@���ԣ��Y1v�?��nKb�D!�������*�T����hˁ+��j���Y\<X7.;%�(�L�bI��
*@G�*Z����A��O�9�׈�K-� �r�o�K�̮.ЕҚ�b밈�#���X�'�@�Լ����$���?n\�%N�RZؘrm.?�.UQ����o%q�9`{�!%�Z`iZ&�l�=�rϱR�m���6Y���t�3���ԥd	>̽p8�O /]����Wb]{��|! f81T�wNl�]A�eQ�%[%�󜢶L�o��t�O��Sd��$ޗME���A��H����̮-�4����gp�MN5�+����Q�?dK阰�`B�k��l���MӁ�:$҂�&i��P�T^�;�x�vr��k�G	����Oj��VL������ݜR��;-	 Ry���faɝ�8���#Tw�V�=
^���������i�k��{.hg�R3�X�f��{2���
�xH�N���A����ˡ�LI��Z�.�h�	~�q�_��J�͠Ґ�����]��{��T�%-V���,'��U���d��{��@�+/�S�)&��y���?�HRa(񕹁�B�5�N��[Ⱦ�ӯ(�3��B����8?����R�D;���ͼk�	������#.�~J�b#ᱦ y	���H�#����I�8�N�~ė$7\�N�9m�qY�oZ>�S(v��CW�(M�غ�g�GS��%�7�
��x��|E{�T�"��f���ˬC�7|T��"Z>8��Y���˙m8��nZ����_���������R�%5������u�@Jj��sX��d�N�RT)=	o\���
�j���݅���U3��;7����	F�y?�J���K���_�d�f��|R���h�$��g�y���p��o4%FY���,ʗ��޻���<��k�k�Ɠ:GX�"���Sʖ�,	#��r~��.�`���� �5o�A�25J��em[ln�I�4����l�����|{���\Ǹi��Ԓ`*��c��:�QS����~�9'b���hӑ,�:�zFA��W^�1�B�����˧�m�t�E>��K���S��cyS��r�ɗ�媡񘊽2�o��
�<G��!G��-�C�wD�*/���bK62iv�/�E<o>��qm���@��v�T{ܢKM��YJ(���Zw�'x����4=�/:�<0�q�\,��a%Q���.�拀.l�3�����^b݃���m ��{�� ���c_d���~)��Z����w.��S��Ҳ�����3IO�Id���S��q��r�����f~N7��v
�jT��X��Ls紊�t��wuK1�#�'���.�?!
e�1�������;�Q�w���\��H�y��)�񶝽�4���UR?e6w���y4f�E�dH~�ޭ�M@ɬq�4�0R�(#B�3@RFA4�Tm��"i�P�j���h�kM�3���)��S#r tq����E�<�G�<Xހ��E<`��}Ʌb�Y�� ��6s�@��5r]���*8r8x�h�w�j��7�Dҝr�h�i+�i3��]�*�i�&�{<�N�'y�/IX�?�	�	w�>�Ù�9���-w�ϰ|6����_H(W��}9k�A�O��%d�zCdJ]M��!�����"J�w��"5)�U�5ڟ�b�����_�gh�Z�,&JM%M�w��UO�;'Ӧ�T��7|*�9� ;�Y/_��/a��	ƃ��(è�*/������CQQ�1��N2������z�����	uQ"
�����j�G�{_8 ��d`�"\�~���Q։��Zw��\dC�7K�V��=�7or���;7_�WT�o���b�'�����4�G���?a<T�C�|1V�����1\�s��O5�2�qKw�k�)��QNW~�0X���:�T�ym�i�R��:�E,�K�����
^1�B^�AyĮ_VQ�2�t �+�*tWD���Q���sbS�a���E�o�����n-�O@q�	��A�E����G��F�>7���>.ϊ�3j�)�b�&${�V��P�lD1Ǉ�	%��"�dH����J�VIT�_�X'H:����N�Jq仾��e2�*�U)	ӶՐ"�K�S�Vu���3���zwɫ}�� {>lՎt>Į�(2`�6�=���Y�;�Ǜ�!�%Su�e��W��P��Nؑ��9�	�8Ә.��|��Ld
F@r:ط5�T��xD��Y�����C����q��}煮+��XΝ��?�4���z}M����K�G�v�ʗZ|�Qz�lWCÉ:��	L�	|�G��7���_(��f|�9!
 �.4a�X�U����S�*Hޗ���q֬z�n����m�p��AH��xD����R?��fF��l��{�yȁ���ͻ�t��	Fھ�
��
2
#12��TU<ha�O Qف�.no0i�e=_ �}�e���]���f��AR~BߦN��{']��U�bHV�;v�1�g���RU͊~çx�{���>�6f�qr�V���i�B�D��(�1�G�P]��8�^J����=f,·.�zTX.���_�Is�4�%�������΄TGY�P�D%6�a��Z���Ő�Tˇ�����9 �y�dbʹ�d/�d�Q���pM+�E���Z�4�=�E�/VJ�[	����ܬ͡$�=₤���>��:w&d�yP/𯙪�ٝ���$CM�q�s����G_ �{�8�0���͌��I�P� P��i<�6oj~�;Z��%����w�e�iou�Q���dE��I�[lJ⌙|ۦ\���j�$�����{e�9�H��𚋷� � ��mpMf"N�Vr(�����>�>@�6�m���&�ɾ���K�X+�Q��5m��G+q�g4�TY{�cY�1��4���8\\�fb�)�~`R:̹D�A�n����d��3�m>��q�I(�V���?4��1��
 �m����'Ċֳiy�e薹u�=���u�\xj��D��ߍ���~h�󥱺�'_f�y�(m�yĦ0ܽp>.����n���(����?�4�f/~C��y$U��6��W�`m��͎�h���D��V�,A)y�٣�nC�k,?Lg5 ����7� �p���A�7d{�j�������p�Ў���PF�]-�*���s��-�H|5�>�1��<!ݔ�ϜwA�f��1ڝ*����綿�W(�I?.f޸�c����H�c��7��E͏N@�����"N��������]Vk�k���}˞7/#�WA�k����$��*��%q�-����8 p*��pT�(zB�*kE{�K�o��&.U�P"TLH��������`7S�s�5�h�Ƃ!�06^w��h֖����9������-ԋ�2Snv�r�^��1��:��>�]*7�f�p�=C&�%:؇����$��_�ԯU��s)൅v�g���B���$!�*Q����d��K�0�w|-�\�K^�� ��1TZr=��/ggq�n
k�R�����dA���P��^9"�$H�?�G���a$ �Zt����x�|eo�^z�=z�]*�	ŷ�O�#�q�UZ������ނ���|���th,��Ĺ;���9�?�u�2�i����ᜑ|R�% �<�y����ٜ)�㸙�Ҿ�]�Y-��?8X^)�/��~.�?�F�G1�q�Xq��%�����7�%�h�����t4h��-L�Z���)g
4Ж��z����H��j�2B��l�H�)$���Ѽ�y���<s�x���\��\���}Qa~����xP��cE\s�`jG~�JO�7��5�/,�5�T)m5,/w��GW	YA���A���K>W��嗢�B܀�!B���t ��n<dY<����Iªӥc<�����G��ۓu�9S.K��r[�=h؎�Pҵ�wU�4��58T8�_�-�a(M=8�:E��Y�H=�h6H���[��Rࠚ�s��Y����,�2�t=��f�d�{��,/W�m�7O�
w���M�|v:���g�D|�#�i���a������$f|v�2�`����m6kn��[!�ȗ�����D��'�,�]�h���aS��N̑M>��:��i��@L��#@�)y5'�z�S�����_Q?�qW��MSd�VdP:���R��.��X�ʐ��^
V�IBw���gf6��CO=N�ZiK����A��A��H��}n�K�PҬ;4%��L�N�<��I���LEK �.'�e�Hf^V��v��<ϐ���)����#> ��L]kT�1�:�Ð����^�f�' �(��}G�t��8�����<s�
�0�?�@ɧ���F�3�Fk�h�Tk�����[��r�����R`=����E�y���JM��Ǩ�\���+�2�\c,���F��r)l<���G�v���[4��-!��u�ػ�<�nh�=ێmJ)Ľ�[�bQZ5�γ.͎����U����*�˽DX�Q�[o娳�j������B�����c1�0��ͻ
���-��Ne_!D��<D��KY������^��~��aTO±
 �[�Gn�dP�ծ#0ϦIw[�z��uNf,�
�AY��o�=Ӕ��8I��!�_�-�[���(i��zbl�?Y�u;����9��|����<\3"T\0���~�\��l�j̲�&d+�d��t6�x^qF��/eNM[�����re����_7Hb�L	B5�p��T�kS�N�]��\P�.��I `�/�a��ƴ蘔;�wA���+� ˶�Z(�i#t�p%�|M1g�GA$A�zQ0K!� ��*h�
�`��FZ�L��$F�I���˻ P=��#������g�����TqŖa`{)1�GV��`	�脑��]J!pZ^c��n��Y%���#u�>�sۈ��f��F�w�D��2��f����4�[�Q���H��%��悃zس��2��Ń���h�c���B 􅁑���Y;C�ϑ����..���C~�X�/�G)��QP�	k*�(#��=��V�+�s�J?x����+) ���g)���b!Tȩa{~�J {����7+3y��0�W�Z��Ĕ�f�K���u&9�6��_.����~w
WA��o����j�d��]Λ�Rڹ����'������ퟏ��zE]�M�^��A6�8th�S��?��Sǆ"ᅑ0[,:���ûΦCݴR�C�e��-5u���&��qtnZ��.N�N�N�#�|@�u�y��EX��*�f��	�8i�L�6wv["�F����]�"���G���;BqN^��O��-vt �#D˦�*�I.�[G?-��q���(3 ��5�N�D	�W�d*��|���y��g�,i6L;W9�3����~��~"��o����;�3��dl��[;�
0/�yĘڷ�_5�N��Ǐ0K��+�u�Y�1��X $݇L�-�eE�U_QШ|BT����7k�` ��Tq�'�Ɛ����;Y�v��w%����Ho�!��
/=��1�\?���8�oQ�_���W�P��T�>�H����>3���'�/}X��i�����*�uf
WC�U5t[}�[���c�F�~@���<w `��i�v��jQ7�U@���6�N��U[E7�'td�9�#�'�`!�io��V�C�|'k�?"� ����%����UY���o3�W7H���'�FÌS�D��R��]��Ȉ�4y��M0,d���� �q!��?h� �0���kox����Q�����'�M�-0�[���3*��Ml+}�g��^>8�>��(�KE�hӬ��'u0Ӏ���㾈.�X~KŃ:��ć��?�`=^�\&��QO_���Sy�tjuU�ۗ�k_�8���{Ւ̤�vM�0s�T(P��ڐ
`^C���v�5R��4�n�ƽ*��Y��j�^'��˦���V�o,5�m3�	73KYc}dkC$-Z�uH��i���D!ڐ��u�9vNwsi�l�>ڋ�	iߣ�(���(��
�Q�%�K;�k.�"r��=�,ec����>�R��M�#pD�� |�|�u�t_�s�!R��h�%�]�̝o���9W{�\�;e�ZD;$��B��'�;)�8���`��f�Y�m�M�#I�I�J�J��Ȫ�����\��9�p'|\������8Cӵ���ی��
~aãY"�����(0��U�f�%7�  �g�\r�x0��
a��!ߺ��7?	r%���=�b����^�)���s3�Y��Y&�Y�a<�i�sd�\B�9A�qW>�evXV'�_���[��J��4{_��ğc�U��_�f$�翰�"�`]��8���wK���C�B��Y�S�ys��<ɭ��w���L�Y�p�uR�fB`=_�*��Mx�nG�ؒ�*_1Q��Z_Dǰ� ψ��a��W�
�eb��-�S����;q����A-o��Uf�5�ѧ�ќE�S����� �G'�u%;��^T���x���o�-�Io#f��O�[5l�{��c�Y��+� ����r�y���!���F��֥.�^k'QI�4ǰ����Y#��5�&�ˣ�${��g����'o�Ie$�!�%9��_���z��Mޢޒ�g�C���hc"8 M_��@��6�!�}��!��?�x���ܖD{�@�G�RcP!�*y���%�g�i��Ķ����#Sn��Wm�8�_�`B�0,�?�r B!�0E��S�����t�o&�
�
����`˽>���Eұ���6[K#N@حRSL�9:Gxsk^���ϊ��o�f����w� 3����8�U�Op�p�>�m���#�7�u9�\v�����8���dK�>�?#���U6��"k�����˔ep*R�1��(�HBe�h�]w�qx���� x��X2�k�Kz��/Yu����T����ƕZ��E��^�܈N9�>c �w«��$V���M�3��o�!JՔ��e�<n������*� �.�%T@�+�ë2	��/�	�~�K" ������]���/9]&K��n����?N�����L��5~�8͟�Z�	���ωj�`(�_-o�xN{$��BK�"؁�����;E�H��i�m5��ʩ�5(��N��7P˫Xr�p�f(W���q����[$���3�\�l�ͼI����v���tm���!7�5�ћ��Z;n�3q�h�F�
��[��Y��{ۑٕ�6h�\�zy�G=.ŀ�ۚ��WB���6�-4
>"�p{R�C��I�P|G��i������;4WI�Ɓg��G�VHD?r8Xh�0�9S��j���^����d|̨\��Y�ĵ���EH7̶�N�O!�9pi��I-�{�8�X��ݝ��\�p�6n�c��|F���YSc�yʪ
4����U���URDgg9[�J���E��<iȢ�i$�"�1�ǿ��fҳ�B�۶��L�A��Л|v�^���4tr���f������m��ϻ��
�煭l�8H`'S�\����J���L���&��V���Z���Yk��g��n����=X�C�._D8>��i����_��u�W�>��E�	d:Gl�l�Imj��O�����XT2o 7�ʕA�G��٫ i�'h"$�Cbh�[B�'4&�E���+�ȤL��C}��ۂ/`����]���?Y�W���o�쎏%�GN�NL
n|`��T����1�����)r|'f���H��V������/��"2���8�X���DH-��S�xlc�	���(��kR��<��Tߪ1�|����;��*�$A~��5]��~�y̔��t��CMc���z)vٖ^����f~��r�A����ʬ���9a�e�F�7~�T�To�wk6P~�(��@��c�|��F\��\�S�gMLB��6�b�,��� �w�v�_Z��:R�ã/�M�S	�"d��U�WH�5� I*��@Hil�	���\��F.M����`d^�/���v��܇;�T�����TT��C��Dq�g�*�6?1�*	7?� �*|�,��pE�c�:�4VF -Z+ڕ�,R���8QM��^1�7��AP}u3��K�t&��m��90�scr�g�;�6��^��CVe\w@RYB=d������׳�Ա�;��Z6uz72�Q�����5
J��Q@-* /ж<���Ǽ���)����R'?��H��u�V�@��O7��Q����2��@.�Ǵl��!F��F	:pQe����d<p�Xw9�8�rg&\�_/P	�8��#��,�ɗ�=�Yй)R��"�nۘɼd��Z<>UW�|�h�AG_IK��b>�ވ��$�G{����y�g;r����}�Wנ��JߥDMAK��'W���ַ������ʚ�+Z���(�!QS�U*e/�P�	��܅�*ܦі��<x�����R�2<L}��8���6�~Sx�ol����x%Kr�h��mwa�/��P7�xp���L�����K������#�s��C����qk`e��\윞�C������D�3xL����L!�;_kW>On	&ɪ!Y+��7J���2߼�����7ά��t��~�{,�>���U2`�U���!٥�I���AZ���
]�nѐ��HH݇R�΋�:�	��	k����f�D̍\�Ǩ+#�#I�7V��M�Ή����h^��'����|C�w��!�-
��l`�g��8}`-�,�3LP	�ȇ������9���gr�bg�z���@��yan8
���43�l�w1_r>6hK�KW@)f�L��
�3�$:�B�i�����(YUoO��� �;Z�/6�HkD+�o�k�<zO9t2Y�5���0phz�Qޥ�ퟏb�r��Uުr�-�# �U�i�{�|8D���R6nR�������g�=|����30�o�e�
KZ������hQ�x�%(�{=�$
�tr�I,�k�� �+���VP�W���ct^�e�z�W��ljK�p�@�r/ٖ��,Ox���Q���eՖ'���Y�mS�~]5)#��0G���P_t����Aܐ�ؓu]�iQ�ˏ�ި�wQi�H�W�7}7o���Vڦ���U�.@z�0��I���"?�O��޵ �"H�>�/�=8�cb@	�� q�Z�����X0GރX�0Z�e�_$PLXM�3�/&��M��¹�>,�l�Y(��c��������|'� �hӧ���ѝ��8��|�Q�o���q.�Pu��GiL����D�>~�d����w5��J�<��,��k��'FA��5�Vu�M+4!P��kT\j�����T�ĵ�[�$�0��r����u��*��PM�;��������yh��n���&K+�i�]�4��3G�I�l�_B0,^Ove��P��b�Ӑ�,_��{��krj�h�Y��^J�,�D����P}�����jOߜ���8�`L������@�w9:\J����!�S�^%H�O�Y2�p"��R#�շE@\Ƨ���kA1�l�J�����I"��t�3]5�ۄ}���[��>q�(��W'ʟ���f�
8n^��Y�D���L9�������� �l#�*���`������:�~a.(s����T�̋�]���!��?&&���q��z�vN�:���1F���i�dqD�X�rƤ�~�FW�\>��{��QFL�)a~�.����q�7};ٳ�2���gyE�n��c5Ʉb���	�� �M�������%T� ��@h�kiW٭R�����2VX���^�lM�ִ��J�L-���MNfJ��X�����5}��;;��+]ޗ �H����n�#|j��WhV�̴�P�.,c+�����ǀRgL�ɱ�mV��bQ����T����"QU3������!f2ię���S��=�ɜ��/�dG0X<H�#��E��a�Z9m@����tk�,i�WK}����D~{�Mx�&���6�ʣĴ(gf��z��8+X8��w�Oy$�]���Iۍ��vO��:h+sg�5�:���n�u�g�%\��l�@Wr�u��X�
ı^����}�1�ʳh�X�b�>�|���mŽ"�^�骵��]~�O�b��>�k�$�[��0Fz�Q0�c���p�i�����)����@H�O�~u �{j)�+���@!^�]�C�Ԯq-��y��o��;�W'�au���RF��[�~�>�������կ(���Õ���~1Fڱ�2.Ғ��(�����/�8VPge�W�ӂE�-w����AË���-ӎ��Z�m@�$�G�!�M�zs�E��ڣ+���Y��噺��z��X���DY-��v��Z�s�Z��÷�v��RMru00���-A#�e1f���v�K�Nݖ�»u&���6�=u�1@z�<�ځ�<W$��@3��X�+f�ܸ�2��pf�/6X��T�tc�|�[K����wء~���6h��5W�~��<5l�9"?D�q0 �.�s಄���a�jW� ¥���>��Gq��4:�X��Dq�-w���[p�>B{�RcB#^�ƎK�}PL[���ۄ�6�{|�U����7�&��"bD��\i~u�K���l�0�;������O�����D���O��Q╬��?A�d*�qԖ�%�Q�@3�@�i���e�@���>�l_��{�H��z�q-N+�&������[��l�m��l 5\/
(Av{yl8O��B޶ʗk%[ܾ�8�6�ȱic�SUT�&F$��9��`�?�s#�w�*㰇�0
���.�xW�I��C㎺ul������Պ�����in�X;�6�N��z�d���h���ҹ.E���6j��o��G̯�D�Z�=��rE�bM��l�3۟�?n4����1�N�\KL�3p�9��"Y�@����D��FGh,p�z�?[$Im⴨7P�.���ӯ�	�=6���Dko���g>����c��� ��V����9)�dY;B>�~-��?�$��`A�YjFw�}������F�]��%RP;�3���D�UC�h�vy�v�5hq��tr�� �jl���U5@�©���_J��n�ؿF�7���`�Z~D@�Q������8#��Q���T���q"�L�/?Lcj����/H�B.�e��s.a>�r�bhv�LD�-&��g���WwREA �v� B��Ovs(&�;a3)�7��M�s�KA˒�$�r�Ն�6�US)������uT� ���^�Ni��d!�jw���>�x����#�\Y�I���V-�s�%�ߴ�X� x
�|�`�)s��i���N=��1�'@
�v	�!)A�n���Fm�ˊğҜ5���;��P���<��#,H4�dc	6FE�����/�J&Nhr�G#	��'l��m�쨯!]���Ł��ّ�e���N�.wj��~l& �?^��pʅ��gK-�ӽ����:D���ة'͌�q7��c�J� �~��#����ǩ�B<��Cx�6���rŇ�a�ގ7$��ͬ� ����h�g7���+.�`�O�o[�^z�96���&�6�˅�����8����(��t��`����R��9͢cQ��u+�a�Hru6ϖA�J�|��ҷ�W�K������!��76���yR�O+B|9�\*c�����Xň½�ܲ�Jc���Q�d�)��!�Ƅ���l�����J�E�j�F;�WԎd8&�Nk�%��/��\�����c�Q�*�4ͳLGu0�Rv�uF)i�?�.��n�����D���ڐ�t���@���/Ҏ�8�Ml*�ۄ~�᚞�����r ʡ�+ei27fB�10%@h�L���ro�^�U_� r	"x�I	���Ѫ�ޗg}��@�z��&��ejM���uLV ���@;1)邓zĹYY��W�AYo��j�5��� VG.��q��>�"�E�o���<z}����I�Nr��:�?Q�ˡ����,C����;u��4B[�\�
�h����眠{>خ|oM�l�	�P�W�-����T�0�65�ص	9cC*Js\��>^m���D���Ǹ�|�cd��˂C�M���eo혹.�L�p�fūN�]�5v����@�Ә�/?��/aD�@e��ȲknG��e�J/�		���Y���sa�����ih{弬W��Z	�ty��
�#��]�ہ	�Rҟ6��{���A��93~hO�������F�'���g��0g$��6`�[�<ۛ²`(o��r�G��e�6��Y�X��_ha	Hb���T�f�.6 A��4(�O�2�~�ܐ�wa�=\o�U2o_v�OѲ�'Y������N�fyE�i�w��W���8�� �н��I��I+cqO3�Y�W�s��_́5���x��u��Z���k^AX���s���u�2�7o�@��|3T��#�ӛK<���K쳈�9�OV�-���I/��C^���(D�£���6/�f��xѓ��O_g��og�ff)
뺵������W�<��,�*�=�hZ�j_���f���l~���A�62�u?����C
�@	ӂBV��?������}s�|���0��K�x���t�2��π�s� �$,p\��(������+�D%�kj{M�
��ƒu:�e�%Ñ;H=��������Q�L�'��Ч���;���K
VI�%���v!K%I̞D�pbǷ�(f�&�/RcV�/Aj"���KP'T� ��m�c����յ��b�ն��[/$Z����~��@�Ș
�e�
P�<�tJS���R������՗M��#�]�O$��岏|�-���K�#���C�.$���l�{Ⱦ=٘�<���o ��Xro=%�)���4c�Yq�:H4iV8��a�ܩ��qlIW����Q&�t�e���T�z�}�<��f �%{���o�s"�t6�d���1)�0PEm֦ͪ Z�v�&5.����5�t!�h���v}��.q�;���*ٯ<�e���~j�>��e�h���4�t�s�S��B�X%�+�-����C] �OV��fA���!���[f<N�q�d��*���y���w�vU*���5*�Ǿ"R#~����~��)�t��l���i��������T%�=ֈ]
���B�(��پӲ�Yɼ�zA5��g� ��:���|��ա�Ě�.)~�Ё�V7n?1P�k��>��t�Z��ѵQ��Iv�+�W�7��4�L:.���Zc�J�y�p���2 LA��1��|2/�O���n jd[O��؈�g��1eK>R�=���m5w�}�p'���1Z� ��\6��
��(n��
�(�I���2��h�8�κ�D�W�6e/S[���j�}�w�G��7 -�%��ܮS%�Ib�E�����̱��Y�T[]rF=|p����w����r����K�GS^�VFx�G�ɒ���KD@�����`�HHO
TN	3.t~�E[5����لz�v�����@x+����*ŉ�Rc�^�mCp9���ī�P"�D�^
å���1t����dMeNC☫.�F��]%6��HuY���X���f{�X�`B���U/X����x�����Q:;���Q�ԧH�i���Ȯ7��@�A�EXp,��Ȳ�o�����$7��Y�H�v�o�L[4:�l}8ǔXhOs^sve�/����$'��L�q;�I�ۂ�Ϊ~�����Q��w-�˪}D�p�����p� Źց�ʠk����z�F�uͧ`�ڴ��W�k��Rq4�S��p��O��A��v�!�ǧ��~r�u�E���T;'�n>��,�C i�i]�Y�}��a�R֪k�J�:�R����� >C���	����X! ݼ�8��������d������^):��y�SQ_0�� n��b���˞��RPI�6�_�;Ui��!"F+�Zr�ys@��t��Н4��iM�(�A`U�č�U�U�ް�8a��7�ML;+��}t���>�[�k�s[��l+J"�O�jŉô��be���.{��*q��m�ε��F�Fu�F�u����%��ҏ�|�r�@I�v9��>\��UsS`���_Sx�\�j=��y�P=���]��7l�`*`�=��Df�z)̱<��ɋ�ÜJp���.��YV����<<}��J�:9�ț浧��s�D;�8v�}=V頰.�" J�S�� �Y�R&d~<BU��c�W���� �Hw�[�y�n��̓�^���1Jb�6��׃�Y�b98M����E������5�i�IS�?_T~�g���p`�vW�F��C�#�ٺķ��o {���b��#� ���Ԛ5s��:��jD���#�1�C���Ӭ��� ��: 0������s*������_m�}b�`����Q�Ձ���J�H��W����@�+7D�2:�,���
���=�jU���H�EIK��	ݑ�_��"�yu���B��,{�����L����`�"�����G�ѓ+�;�O�Mg�����;�As�*@�DbV��MHז8���x��/fIr/�zޭ�@qo�~�
��ܸ�)�|����
q���&���N�������v��r}�L�u�C�U�Ј7>u[�PW�OK%����5���e�@�;�h��l���l��,�2���z�S ���꣭�x�|+&�|�&9t�xD?�ԍ{��oWq^'	�BҴ;��k�ۯ�jM`oRE�%��)!�KB<lw%Kh=ꬨo��o+&JN[��zB�y�0����]�m㠄#DQ,̠x}�.��\�&�5cMFx���~� �_��l���9w՚��o�5�/�f"��m&�x;��
���*�Sj$1d:����s�o�)�Ea��\f�����|f`���S?�����*"G3�]=.����< �T�.�/�%VGxW�Z����y�%�e�ZR�h(�dv�?�����پ �?x4�(4`�uvV�6`��W4v� ����e�T��R׼���!��[3h���ΐA��D�x5�g/�������3�8J�|7��$t����T�X����|&�0��$Ϫ��q��Xyq����2�r�����C��f�#՟�Y�\4� y=�؅梹bs��Ѡ}�r�'R\���\�)�;���M�^�����9�xC5<]�fy�?F���͢O� ���pm	�R�n��[�)/�h): )�$q ё\FU��~��u�����C�Ӳ��L]���4�2������C��i�$%��R��@�c�D���wAQ�X�{^z��؜m�Q�ވ���@�i-��;��E��F���X�2��0d���{��#+��o�I����<��d L�6o���S���	.���*5��3��
S�L/vb�w����%Ĥ�S�����{&j�ByUT�@Z�"�����"��2^��c$���w.�4�nw5�l�&�XRv�x�v��{�����/�VNT� �z�'p�
�k ���\�t��.��P���]�RL}��0��[� �"�?�z��(��� ]���x҇vo�~-֬j�n��q��9t�;����3�� �'J�q�$)n�oڵ�b��w���PI3��U�.*x�E��#�_��N4.�OP���#�Gm` �}�+�"��Y���<��C�7����6��?#�p��1:yhsF>s�(/��J��G�� � ���+�Y)/��!��-�n�����g�zb�p�o���@Y���5�"���1zpl��L�C���h�S�H},an�h}�	�X�m��Q8I�s��k&������{à�F.
}ڛ7����U7)>ݼR�e��'ӭ��'�ϓ���j�#BO4�l�ZK677Y@D�[xN\���lgV�[;�����p?�{�����XR�~��)徍װ�-]���߯1&u8:#�s����:���o�0�l���r�.	+Ў�d4H��S*�R���,�|��!e`^��*φ겗�a���AjE�\4۟f�#��2����7o�FKެ���p�d���-=.�JoB�)�f�F0 b9w�g��ڱ,E�C.��Q.ҽ�ѿ�yQ��	t�<KU�*�m#���M�լ����yL�-��X9�Z2�N(��'Z"2�n��)
��x�)̿���F&�gKrg�Lp;���Xg��b����%��?^Ҫ�i�L�}Sd��bJ�5D{KNE?r[���)-q\!�!N����p�������@���6ud#���4%&需`F�kx���~�l�-�Э{��D_�+6��"eYr�pI��M������f��\�3��s�PI��Qϑ�UF��q	>8��b��	�l8�-ؠ�>u, zc56Q�m���<�c$�L�i�%����{e-��5�-�l'��%�g�l�(v|W�V�
=�����?[�{Ck'�7�&Nޛ���taq'6'�ҋ[��]�q�5l�?ʞ<+>t����4Y��>dȓ�.�X�l��	7d����7R������);/���G-��J��׮ᡃ�5�@wOu�TXo��΢?�$aũ��T��e�`���y��\���(�I�+�����}�jv85Z�?���F2�t�[W��~\��e.]�J��h�°�G��AK����.��� D����|���]��~Д�2�<��}b���ֹ�|~��_�lL�k�*���!MD2Cl�h����H�U�Q;io�N	.V5'|Ԕ5��]K���J'L2��$�Yg��M����1\�ro[%UnB�,��`u�^ϒ�B�:*D��k ��V���4:�M���N�2�E[ k�QۮḲ���<�<�
S�HcnmY�E�[�Z���'�˱�y ��IcJOv`���~�]��f��ϗO0,K�Ħ�ANbfZ�/���}k�(��򔈓�NĮ)�5��Ai�l[��s�@���7�B�v=f$^ATe��\H�����(8���ѳ����|�ػ�䲒�ŉ��1����q��2���,�i-:�3Z�Ǳ���=N(��^Zt�@���sxCv�*/�\�y������Pª.-������
��Ӽ{犥R�����WE������0g�B^MV����]HG?K��7"�؞�-/u?ʤC��Z$��0����]���2y�b��1��<�ǟ�Z�������s���隆�!Z�t3g��chNi�.����`�
T#N���~�Q��� Y\�nzʠ�PGN����Ȑ��!Sj0a2�_&^�]|����BQb�F�-��^j��~e&Ӱ���YG���_2-���K��	F�[? ]ĂZ�[����T�a�,#���hu[(��}�������#/�1�$:	������C�aJ��-[���u+���g��S wg��g��; j~�&6��.d&�(�/��-�O)���	�l���4�� ��MaL�ʸ��(�Yjh�g�A�N{�A�{M�5����w��nM�DG�G;�������
8;Q`R��<���V����o�����(�u��2�c|=oo��$nZ�]��8s���>�=(��+F�$Fй'���ҭ���|hJB�ͷ�OZ�#!�����bCP�R�s��J�
�N��@Y�f�L��_[��s{�{H)o�"Ws���}҃Y�2����F�)b��`��W�x�F?.�+�6ZDN,%�Hβ��A�Ra��q�"��D�X^g2M1l+^BK���M״��Cc�c��:s�G���q�mh�/����Yk�N����+柖͇��,�3�4��G;��'x�3?�
[
GZ����rg�ͻ�����SE�{�6i2J��]��� �tU�Su��w��K7��8O�1��QXZ�c��Є mpi���(K{AVԟ��R2��}6>ˎ^�<g��5]�ť�&���Rei2���h�
�uYaU'8�/q)B]g1��$Lq=a�%�����|�R�2J�i�x&
¬����=��x�^�V���6��}%0�����0[:�[��'!N@4_��3ʊKbס��N�\�_���c:��NZ�+Z�g����bu9h� ��m|�'F����XRΣ����8M"|��#�Q�yʇ2�N���g8f���!p�˝�/1#*j(a=��9e&�bb(�3�|b���K	�Q��"ዧ�P�3���`Gn��b�̈́n&&W`o� �d��+&i��+��/Ý_/�?���G�;97�S��f�n1q��W� ��+4.��4ja�"��B�w�x�^وK'�Ӳ���7�eJ�Xʘ���l��)�ؘ��,C^��O�@��֥�q�qhf��!�i��Nኀ�����xl'�y�J���(��e`�|E��ī�j���Q�֜W���R���f�~j.�L�ns|,B�<Ā_��c3�=q�Q��i��V�XR�>둽l�/�r�}_FJ�ƣ�k@����ɘ@ �$��8!��}nZ���rhMN�Qg�}����[�`�R�s�YGZlu�=��a�X�R���w�J�W���IVm�C�����p9zw ֻs>�e�&z���o��jRWz������8� � �~AV�td�N�p��0�x7��`���g,��1�r-�fb$����MK����EMi7T����KN@kdꘀ�jMt����ܢӌKk*��ʘ�z=��f�����F����/j�4�%(��>�^ܠR��.ޟݶ��π��G�4�U�q-n�C���e!� O~E��z]��P���jasꣃxB�R$��f��>0}k�j~G�F�25 �M3@3�3��R�-F����q�"K��{��,�&��3g�M�����E`�l��-}�s��2�1޲�&�.xM���U�ٴ0᫧A�K�Z�1;J���NÃ�7���Vp ��9����0(��V*�£1�G��}Jc���ˏV�[Pp�7��H��&���h 1�-{��F�@�ի��*M�Eq�'��%�>?m8��WU����X4Y��k{�ĉi�)��VS�FjҨ������CͻOcu����IY&��-�����w�K�2)�9���C����f���2(��n�!!��Ǥٺ��u�p�L��t�L��i��8t�t�8Lo9�?;s�+9�ZN����`�\�l�U�.���]�������$h�l3�ՙ�4� z�!�ڊ�6�r1}η��4
����Ω �*����h�r.n���T�t��͵���"����N2Re�	0����0�Y�فؼ��@�@��,�<�	�t LG�W��=�� ��ۻVW�Y!�X�((�Z�e \\:ǆ�u��L���9���8�#��7����&�����|��@i��t�����DÕ��F]����$��H��8V&\�n��7CRf��gD%$.B�G�`y�0���Ξk C�aC@af�~;k���r��d��.�9�B=$t� m�y>�'<�w����,kQ�i��_���X��L�,V�P0y�>���[n�oد�����N�믂��]ȋrXR��zN��֭��tޜH9]�����'+���Y�*�x|X#��{o�Z�\���M���dcr�GÿP�
o �#�^3W=)J�X>���O����t�$c��<�yͳ�Y���z�F��C#��)��^g!�Ճ�C�?P=�.,�Ε8Q%%�*�46�\�#�)*ґ��Uh�%if�`5~�ݢ��.��!�C�Y	�$
�I �wrbЧ�(/�k
������w
�����'jz���t^�S3���w�s� b���Z�r:����U0#��z��b� ��Ùǭ�Q:��h}���d�w������o0�����fD8�Ŀ{?�yY�q#�A�0ly ��fq|��I�VGB��Cm���~a�ox%�!���� I���[*��5�L~���ߋD��X��J]�M���d�o��ݕ�8�53�+8�"��)�]i�O����>I4��'W���U�Ud�X��@� y󯹾�
O GN&��]��lI�曑j�Q36˿�����0I��y�64.c�4��Q}޶\ 8&D�#I31�^6ݘ5l]�)��1>����/���S����x�r�GJ�
�e�W6��0{�Pٔ+�c�3�-��{,MO�������^&�
_���Y��Q�Ԑ��~�}]��N�ӊó�0��Ht�����5�>���v(��Le�=�N���Q�����t�[�
�H�G0��C��Sb�+y��H�tr��p%�s�*7GA�.�����Ui�2^�[��hU�S�m����Vv*���r[Gѧ"I����l������Q�h!�����|����!K���OAng�;D(W��<���a�Y8�+��E%��Z��؁Y}��K��j?U�9�Ψ�66n:��&N�h&��Ӱ0��zaQs9=�62�QT���/)�ڮ�.3m�PH�n}s}&	�h�<����W���ew��}�H���,�ZL�rt/'����E4���5.��*�^0��q��S�[��q��1��g��〻ٓW�)\�m���{)Ǯ���R&YJ����/e��>7K��Yx�Q@�ܫ��66��ˌ���㠛�f�����կeV���%v�$%K�︽��}Ɲ��d��g�&E%�TҞ�%5 d�Q$�����T�wZ�ODfj�7��d?)L�dys�>S���t�����$�ތ�I�w"��bz��N3Ba7D�\������ %�:�L�����@��"izh�ӓ{vk����2� �����z���bU�W�#Eg���X@VmIe3�K��r����tR��U>�<n��ݫ�5vrVՖ���,X�d{��s�[��gc�r���Q�*A��b�X7��3����t����K9q��N��R�M G�8h"9�;X����F9t�"�$��.�V�P,wkMم�:�t5�gwp@�sG6@c���S��` �R�y��i�|�|���Ib��;uR-��
���1��ih���?Gh�+dCf����2�$mPk0]�`�l��� ���`������4
��K~�h���k̽lw�Ԇ�$���K�M�v�^��='̘x*�R_�{)�5�OwН�����M��R -:ұ��z[��
&�e�u��D��H�q1>	���ӥ�(�d�2&-F@X��ʬ\'��U|�qmਚ�N�[�ۥ����0^+oc�(����g��1��1 ܺ/ΖE��^@=)���u���\AQjc�M�ɨޛ�_e1�E�������O:2��O��-�P�\�^(��o�Qv2:��k�$F�5���0��yl�Gc�5��֒��E�ӻAi���� ;EJ8Ꮌ"ĤZ�%F��M�(�m�.���¢&>z}Q�X�Ě�q�D�j�}5D�W����A�� ֬qB��WΧ�l{5h���L����8J,ס}���P�B&^��`�*�LVy�n�4��xZ���1\��#�+*�����2��]��.�nS�Ȕ�	��M�Y�S���_N�S���_掮��vD�)����S�C
|�����(	ە�k!*w. La�oX�w�K�[B\�r���e��csL��F]�nil�@��>h㡻�t��%�w�Q��Nb)|�(���pۀ��tS�Cb٩�[3�l��Q�&�9���r�-�(
�s��@
���
���p�d6-�����wBт$s�+"O�5Z4k�s�H����PUb�d�9&I�5R��,>�����T�ʢho9�ElR�Q^l
��:)��v0�^s���OuZ�6/`�&ͤ����ɩ7�$�5�̣����_��VdtC�D�y������6��ud���԰�V %�����[e��e.�2[޿W��m>���Œ���W�7%�A�$1.䉵l<	�S�U��k2u�25囌�|���u1��_3��x�Hh����6�X��(tэ�zVD}ߓ�sY���Y`PSkҳ4���_Z��
�Cx�Ļ{`����ze~��������{Pv�i��f0t6*��O�p5�Yv��Qi��P�ЃF���~5���y��
�w�(�4�
�C���5�8s�Aj�t����w��51o�\�����="��܋A'ID�F��,<�m �l_�x*�H��ӚڸX���� �[Gc�W�@�&t��'�����������"�O�՝C�Уs�%.�ű%���A�
�H����5��-��'3�I�����W,P#T/������o%���a�ĭ���������%D�g�ݩ���b ��91(����l B��
l:�m�c�yKJ�X ����������D\�r�[��z�A�^�p�R݃��B<#k^�O�ސY�#��_���� �NŮ6��Z>���ri'8�ed��?cޅ��Y]
�\4k0�	��f�z>�Y9�cm4�_��rQ�[LoA�� Y����m���C����h.���>R;��A�>� �-'Z��d��
�pя��%��ʸ��6I��0������|_Y�ӞK$�'�T�A��� կ%\���v%Rxvɨ߁����������)s�/���ٕ�8�*��#��L���2���p'	8}�۩XiY�6�l73��'"Ӌ;s�I��0UӖ�h,{��@�:w��Q�+�D�������`v�����
o�Ն_A��i�]WtN�j�F�ܬ�Jz��% �4�)��yK��O�o.0ݤࣵ;
v��W	*��X.�>uU��?e��ҋ�o��"�J{sN�B���=F%n��g�t����ߟ�0����پ�b3dz\�/_�:�@9�%g��#�2�?�_�?��k!I���MP���9fv@�X X�$�s�[0��V!���qv+��/��c8R`��@g���ZZ�h1�w�'�P����V��|~t��Oa�:�G�!��1��qB�,����*��X�|�@�p��#�;��&�;	@Y�OjڞX7�����W$��>`@���������P���P��S�q"�v�$����A�'��ì������#�:.��Q�u�W̞_�X<��_G�h����h�~eM����NAY;2%]z�Ϲ8�k,���VF���W�q��Q��x�\�4Mb�ʻ�	�3����T2º��ށ�ˆ�j	G�x�3>�6��U� ��E�ǣ:B�ׯ�>םf[�W�����E� E%u�a��&��j��E{�
~�6��¥��ag����'���w_�����r�R�����C��s��y�G\�FꡂC͟�A����SV�T���6�mn��y�7	��pH;��-0)��υ	F����O��x��.�d��s�ɏ�E.��L �2~��bI�l�#�~�v���>�nĊ�`�e�&c�����\1}x���x�8��=��t��
rx*�ؤ3�������41���)W�M�׬@ט��w}h�ˀ���Ѳv����#ѥ��(uw�c<���q��^\N:����!^�t��؎nלǃ\2jl�c�.\|��8n�ܔ��c�E�o�����(���1��#��J�˺�|7� $����׹ �[N�"�ݦl��*� �wU��x��R����'���e�%>�PNI?a��ǺT����؊ǒ��������F���>��^-��uI2�u�z��H�x�`Ӥ9���Q�HN�����k:}�����q%}V�$�l�H�� 8p��a4L�8����:z��ɵ�0�:R4���5�g�Vv&���SqE1��N��O�����UYbs��o�����j<K����{�Z&N4C���)y��EG'b�Y�����2`�O�LU�4�7���Z�
R[H/D��آt?�ˊ�
�}6�e(��(6��>Q���,nބ����S1� �m�S-��I�����S���n'��aT��Š��0<8�]H��y`�o::�:��?ș<pA�p�Q��! +Ri��X8Z��:�g�-�~L�, <�r9B[ղ{���M��IY-����ty1�#k�W&��O���E=��w)��fC��`+��D�����v~w�Η�<���&���y�H֫�oT>ϧ�(�*���S���"5�Up|	�o�z���)?�t�u^V���]�n�X<�6`0E
�n�W\.E�&�l��~
�kQ꛲��5#N(�;�=!�pz[b��EƉ��x���E<A�U!:��{0g��7 �)�K�_�;a����6 �(~g�%����\@c����~���`}�h�{��Ne����ǽ�|��P�\�SZ�\��e�rI��xu�T��PB-��Bŭ�Ji; ��ɍ�śn�5�`�0Q�� 2ɖ�:�Ԏ~�H6�1���#�|��^f\8�r7RbO/Ǌ�Z��֒,6�����F�f%�}1������W���)_PhGd�tИ�]�g?��e 12�7�2h\���o�_��߳�~����d�(i���3��C\P5N���)� B�QyS	>�AG?[3H�!U����VQ�5Ƥq3�`��o.�v4Ͽ�K*��䕜hw�5�`b	v�����g0�����L����=Yޢj�K���`��J�c,��KO��Xuo �|6��H�d�X�=��N!��)��&�_i.�_1aq�Q�v�֌APM|�ݬn�Pʏx}}��f���ܦ�c�O�,��l>k�ބF.QGR6�3�:j��bpo�}9��h2��'�32�`���3ʈ�,{��Luǥc�����0��Mᑹz�㋳��!��Xr�n�O �X�qZ�B.�*��D`�c����H��y�_��NX�*��fͯU�&v�uK]�c�4���Nɒ]ЮF-i� � V<�����e�a���`X Z�?���xm�y���@�hLWg�h���6�����)�/���	��2�
Pp������v�2
!Q��'n)m��Oh���|��R#���C�<s|��/�~�(�;~�$B�I�n����K�Dѽ�q]��i!�m�YJ�g+�|�QH�]�]Qծ�ңT /�~�j!s������d!�.KdA��J���ri�8C\9�c�.�:/@�ԯN�=Zlmܼ��\!����nO��'i�>��}���#����
�M��pO��L��X������2�E��y糀�=łF1�}M�j��t�4ŏM� ����}������?v1o+,4�!�ʃD���)'���y{>��1Ȕ�Xu�,�Y��-h�6E3��}�f���q�N��^�5�vHg����]��d��+�f�IG7�ۥ�� ����2��V���ғucM�WA?n���?��c!�H
��z��7Q��� ��.������l�d�A9JNM#��$��	D�3"HHfA�(a1m�D�`-�M�P��3[���jZ���������v��&'KT���v��$�ݪ��3`m7m��emO��ረ�v������`���T�[�$�@FܩV����!/����ǥ�7�ۥ���)��3F�P迸z��ఉ��@�u�T�)��5�̺�9���t�w�b�q%Ǣ�7
q�꩚$\X��� �FsZ0s���(g�����˛������_:��j�"lJ3!��>�?�x4��@���DfR���_��e-��h���Z��&�Ӽ�`焆�4��Է�xj����z��j	6aK�A�e��G�� j-��]v(C�$V�.��yAv�B1�X0��?*0�$S,9���VN�=�B4��Th�h1WH���kĸ�5/4��+Z@*8�6e�Wu0���+8����%����ofo�B���*�+~�W�`����e~ڻ�����f�j!�9�Axߣi!�%��'U�[2�g� bE��"����G�_�>-�n0��P��hۺ�Z�����h4��HW��͋�g�%��+
�����a��Y�ka���Bs�EM�.)?��;�Fb�HS5�g���΍L�f�[s!Y�����$�Xm&�er����0����o;B��j�R.�'�U����RG�4����S~�ݯ6�K����K�;���gW�6K'��^`�������k Hn%�N��B�S5A���858�Q�i����G֟,���"�9�	w�ڴ�N.��;�Q#�qZ��p�'Ma��ؙ���X�M1��2�1d�Ѻr�,��	�OvΞ�����<x���U�QL����=���8���?˾+|4-`\T�b�@��An1W�Y��I;��A�q�gSR�&M[r����L|uª�W��kW�L\�.�ʄ�B��	���o)Er�� +R�B�
 f�ѿ�h�5��M}������bڊ%fޮר8��^���˶�څ�UA���H�![�4�[����<��U&O�m�А���9ڟF���::�㖶�����Pȩ���m�n)�ca����g��5G����KSR��-#�`q�O����3H�!�S�S�p�8�@��+i��-��*��KC�U:���Z4�sIBYmBy��cEk�U�l_���'���,I��ۋ5m�Ÿ�qmL����D����y��|��dnNR�Ɨ�4
�B	�����B�B��G�!f�W}���PX u�un��{lM��$�G�)��G��u��{�R���P�T� jh�)��|�\��cg6�|hdL�����z~E��K9�u'ǎ�5���׆]��r�.ÚI�1�fo�����`�1��Лѷ��hTȕ��p����$���7�$����Qj��/<�?:G����Z��r;�.b�Ug:/ E9T�.�#A�k�� ��$ E����.�����&Q��2�$�F�|�D���T�z�&�,&�.�HY�{���G�}��#q�]��6}����7eX�^~Z��o�Ѩ0��5��h�=GvQ�n��G��_Y}�Zn~+��Zy�.�kڰ��B��jK�I�BD�n���	R�1�J��4�N�t̅���yĔ:ac/�O�M0c#ۄ��=�}"�߫�*vWFo2	�)����W9 �]Y^�9*����t�˛��~̓��P��x�Z�?٤9��r����M�_̰	)�X9�l���F�2z�������[­�l��(z,�,��V���겚*��i1r�h\�.��բ�<=����'~�VD(�_?<e��p�Տg�� ×��';|��\��I�o���
���0��K�%��3� �wV��J����\��	�$���~���_�«����3NF�i
��-Ⱥ���<z&u
<�c�gr��w�D%���������cb�b�4k�t�s��_�=��8���[���,P'/q2\�z4]֝0�Uo(��~
�.hP����S�=�����k�0�?�hh4z�p�Z�O}yO�?���~������'���H�J�Q�c1~mQ�p�� N5�B��>'匦w�S�>���/"%W��+�):y �(�L�nv�X�AF%���e]o+�*��q3���� :��e��U�v>:ڙ���&�|��~���D�-z�45�
�sO_�w�k���\q�`wxل��t�f�8N�C���Џ�kn�r��Q����Gl̂5��kE�s�����g��;=�{�"Gl��IeۦI�L�b��r"��D��Y�B^]��yq3���(�Ҏ:�dj���(i6�B񜔹O0���*X��}�������Hv���v���.l�F{B���CG+z:���6��2V��f�rpJb�]Q�I,j�ʀm!�[Б?� �BÌ�����ۉ�mR�n1��Rd4V��.�CF��?8��fQ�@��� �CLf�V��|�]0����4z����f�����̑�ܥ��b](c�����cl�4E�*.�|���U �`zI��ߖf������= �*�D�ౡ�|���A���ǣ/=�Ž.x2�fbЍ�҈����hKl�5C�ݟрp�a6��N��l�����+2��K�I�K����8ƚ��EX�����B�ɰ��G������q�3˹ϣ��"�W�V^�������n�]���=̜���P*xE�\�?\y?�A�ld�0&�x)���5og�7'�hD
�HJ�e��b���,_�Ƌ�FW���sp^�P@�j��~i}�|����!��-(֋��{����p�2�q����O��`�ד�
|x�'m=_�6�D]Jx�e��čH���1Hd�!p��JbAoQ���O��[(!.�G�ن�!�J�BP��zTơ6��-4b�O/��X#���{�j��n<��T;���'����+�H�3��#�������۞��������@'��O��	w�D�qz����/�G���b!�;�Qy��Jcz<�	�������W "G|�~vQBˁ݋�Ic:t�ᩢ+������`S;-ڿ3���v����o��Q���쬃,��`�j�N��'R	(v�#U|���A+��t����xHBqm��%X"�����*	�K�Ŕq��뚚h� zDʜU%*�� �$�x�U	y24~La��e>QmIo_��E����/TC�砑�ī&���T�TX�6z���t(��͛�� :�� �D�it��'o��{XB�hd��U�Vn�M{<�̈_�����^���^_'�����%}f�R�sl���/�J-�H<��<$���p��
C�9��^��E���.L��nʒ�V�.&��,E=�<��Z��T}����S���M�>�Hx�[�g�~�	C1h��I9IN��V�{�P(�Dw~}�._�ۋ��d��@�^5�j/?�\&��l�;����#q���/��L�Fv=�O�k���b�KZC� �u��%|ˆ�T�T1�H�}�ӵ9B;�I
�ܟ�έ�]Q���R���Y֢oa�	_\���*�!�˶i�� }�'�c2M�e�Mɂ��C�ٗ����,�ɘͼ�}�W���Mؔtǥ���]���0��fn����\���Os!g�Xt�!��o��xe�K��+� A�����B�ÿl�D��'�� ��S�D�[c��Y��1��]Mw�#�?�[x�o�1��J���e�L�JTy�L�'�/��u],a�#��E,&���Nn�s��2��������,�2�PZv���}���S[V3��S~g�#+Cȣh��:2x{��^/�:h��v�+���V�}�[j���>jḒ~˧�������D�̋gm´�c4�n|�[���6ڿە��T=2��z���xlM?�g��e���U=�#��5�|�Ɔ@�N��(^4km���Au����ڕ�)= qS���-�"{�B�
�u�"O7��a
�����İo�57}hyj���i3w(p�����`f�J��:5�̡���]!@�m�Bc�G���$5��ib{)S����JJ	q���W%,��h�鞲��� ����>����o�
%��&�5�yҁ�� !햋��Cݣ�!N�F�e�"(���<Y�D(f^�s�������z{`?�O�E�lC�d�X�p{�3M8�0\f���P�j�{� j.j�'���k����q��o�+&�r�6��`A]��\�Ӏ�r�
K�w�t���0Hg���=�?�V��R�1�Ľ�����<k�a��J�![k�~.���
&b Vdu�qwG>�(�7��6�i&X�7�ˈ�%�a�1(� �@m4��	�?��=�����d�匥�v�}c����9"؜�QԽ5'�j�ߐd�9���%C,d�jE(m��T�	��3	Ӫϵ.QgV��6�E\�72����P�zI�U��t�X�1'[��ˈM�r�":�Ӈ�t�ߑ2}2�_�;��*�3�,��FB�s޵`d�F_3�B����up�\͔�D[9[�(���^ƅ��}G��
�'�?3�"�[
3���e ��:\#��UMk��d���ϟ[T���sTF �Ʉ,��Er����7�/~TF�gR�X֬3z��4��s��9�^�xj�̲����O��e:ĥ�Ac�`�܉�.��ֲ0�Db����e�ӫN�:9.ՠ�7�� �{q�I�+_߉7�.o��@敼}ZFuZ���,�$Er��	d _��f[�P����$�\4�'�J�^ٓ��8�.4�]��/��0HP�mM9y��6�^R�^�<��R�4�F��E]����+��]]
\v���0���a"8��̱N&��,��y�,��	d�V���~%c�듚"�����zK�l�wR ��Q&������+���%=���~�,��T5S�܅e���oT��V�5�s���j�����~�c$r��nY�y<A��	K����R�����*�}��G�����º�ާ��a�[���3
{e��D�X�e�7�E	
������\����:*��'�cb��M�~�Œ�{8�~�y��}�A
����pT8ʿ�����-_��C{DA$3����)�����2��3�#���?~�"�8}�B����AĻ��������,7'i"�x��m�W�alM��GU�9)!>�gO+�y /+�l]V�iӯ��~Mr	n}i/S �!(¬���$E>c��e����@ ����&V�6e�U2�}��bM��L�mO{ 6Ͽ���O�@�܌̥)�Ę~����öO��BD<ih�|�w�=����V�����@Y�Ρɒ����~�z����3�)E�z���|A���m�heE���h(�H\X���(�^���d���ZK瑷f�W�b/�96�e��^b�K�����=�6N��<V�ߒ�GnҨŨ*�?i�;�l^Mj�ɼl��
Sy�O.�� ����_�&�q�W9PT5c�+F:��Q��YaB*SO{H��h��j��mH��S5;z���e�5�'�c��ail�
⚡��}�z�H8��6dz*���ɪN�z`ω�C�5��9�"qE��Z���Gre��-&�v'�
���m�
A~F_�n�T b�f��VXa� ��A�uL%	�O����X�B�C��6��k��3����at����`�V@��]?
�ʲ��%>���@��g7)�]2�-��l���zs4�1�?7����[���P�e�vx�B������<Z����-�Z�cy]N�|=�B���db{�h�s�Q[�hI�.��G�g���H��S����[�b�씜��?�߅��4�꧔-���H��ނ��z�U�#w!
a6��(���7��4�D��,�G`�H��clx��r1����j�9K���*�I���3��pғ��ߡw �*��?��Ԡp���h%ڧ���N�k��+C5���c�a�
5�������_jq��Y�"�.�1S��ãE=Q@y>r�����l��M!G��^�~��I1nN���F^ ��,�޷�L�Fc��*?q\�n�q�Xt�ɘ������TDŜ�l�����{����SE�i1�1S*~�\SViF+��f���n��Cښs� d�ؤ�FÓ����J@�Ո�Ђl���~F�7��,V��F�%���f��Y���tA<���V��6&#U�Af�G %�]�>8t�S�j��j��2|�v��[|C���K�����L��D|.�~�w�HqEbr�ַBv�0!���nZ�ب�iUw8ׁ@�ԕ�Z�Z3��o�wt��ن�H�ZwK{���Z���Т+��7B}!�ޠ���܊J�����E��{@�+'�ha/X�r�]=؇����v�-�2i���	2O�5����2��'u�͠�a=���D'dU��Aeb��BZ���T�i4�]@<�q��T�M����!ؿWk[�'��I��c�H��w�w�%+U��D�Y�k�D�<���_�E��SYR����!{Ь�>���>n�[�hf�8�i���ٙu�v`F`2���:6���a'C�z�&H����̇�L�''S�x;
�P<���2L��ϴ@S���:�2����3�>���ds��d7�Ib��۠d��$Ǘ	o��l���cUK�WW����dށ�W8�� �J�A�4ueI?����:1>u��ݺ��wX�up��}�����̏5�+���J���Ԙ�����tV����
�4?����4��IN��T � �=u�5�/���o2_���H	��Z�å�}�n����q��wc�b9Ӽ�TZ0�+akrYP�Vx�e'� �����}����裾��@�n�*�It\�I*�@S���2�q��'ʲH�&,�RwhGLJ�Y��T&�����^��V%�F�y�k?i�yB�;��E��yA��f���c�kpFd ���W;����M嚷\y�������[�X������ƣ���u��l���弿v����0Ɨ̃+q��	S���I���5�r%
�D_�G2֦��4�/k�&�Ѳ{Ԉx�:"�=<�O�r���S���vw�0��8�PQ냴�1p�&9'#���e#H�cj��G�c����M.j������繫G��_r<��ΰ�Q�35�@Z�<_�|�i�]�~L�1����|C �M�L@u�I۵�Q�&���D��Q�W��h�­��e$���>H4��!n���^���jtNP��K4eϏD�n�]��%O�uUl��wf�S�2kϰf�eo�u�<j�|�t������R��(�\�X�5��*��3E��ǣ�w!���H��y1^~��]zCh�b�l[�����t1�Tݞ�4Pkln�4uZKJx��b����vҟŽ�_��v�>F�I�C�a��#�@F=��f��4\D�mw��t/��[g��k�,�7F�[&P!��:2g0Y}St[�l�Z�W�0c�]|���D�SQ{��~|y�97�j��֦5��;���6C�4)l�`$�0���H��դ��2y�6��k
e%��WE��lQ�@E�m~mp�l%��͹z��p����� ;�C��>4cmӞ~ɣܣ����MqD��h�������Xj`
H�JX�f!��%N#�2
@r���^�4f��^���'QV�rju����Ɵ�Gܔ�gZ���[�|7�E��v�oi��Z=Ml��9�����,k��+�d���g�=qț�ڇ<r�����p~c����m��2�$_��r��s��Q���x%t(��g�����hw������J!�{X�7��I�2���[N	��:�G���KjU�C}뢐�Ο�HF���	������� a�ń*$��oH���G	y�z���U���ր+,۸�̃t��S.�u�GO8az����@]Q���a#V�&u�2�ݩjyX$�yV�!1��LQ����8���kƤ��(��gO��!�.��RWI'���˅p�����c`ũ��y��m���&�e��A:^�`;�����&���>��9{J)f�3��ϢXG�ƣEo��+~��Y$(5n���P�n�46MĈ����05Ia�+����5��[�h�[V��I7*+[YǍT�i���:�d�ݴ/9��X	tXU��n��Q�&�,�.{ /�
0&��B10=X3n�c�i���}8���b���i��wePr�Pu�_��G��N�w^���㕂Y�`j?�/��l"���|�L2ű�l��"z?�?ʮ�=5���l�F	YD�G��H����Jb-�B�/1�G*�gA6n
�bhŪfW��M����9K<��(ܢ�;���s*��#	9��)&�ڋv"���G��}����/� �残T�?~I�&B:�*<x�F[�!��^1:��[P�MP;��X��*��6.Q�°Zs�e�
�!���٣�;��hd6��z?�����p�)�g�I�9�T�������}��oG}�Qpb��'��::�1\����A���#*i�t�����"j�$�N�f��*���3)>�1�-�~Ma�|p�`��1��fS�.�Y���aɅ�L3U+����8�ZO���ـ��n'��Q�ܒWyf:��8�M�U�ӓ�-/5� �{줱�a	-�xU��Zn��a���Q4�:5��u䋏�IW!�,9q������g�2OI�@��V�S� l�/���<�x�I�ˉ�ޣ[hcNPf��%�D�J5w �|��m��#؎�N��I7(c+(")��SOx��w��>��_`�P`QbC����	:�2�Z�� �K@����H�U[+��]q�']��_�Km<�����������۸��I���W�J�6(�G�q���\Kn	��o�i����ez5��t�i�8�T�_RQ�T ��J�O�U)�)���R�&������c��=��\'*)~%�K��R��
��ץQ��鰚;>�r����.TL^֐�<F���zӸ�����1	��`]�~�MP�[�b�� �P8!�Xz��Ί���z4_�P͕�|��p��(%�I��']�u� ȃ��<Ņ.֔�3�*qt�p�ADܒ�d�a�F��l�GsCYd�V�o�4l�H�|��1���L�%2*\��iT%��&�@[|weTOT�C�t�Dq��uF6M��A�V:@�y2�߃�f.���� 1�&3������S|v�����l��롊�ׁ�X�'�頧Ѹ\)öξ.˲/5���@>��?�hoT�^�b��La���uFcz���*&F$W��a-L�������\����{��6���2��Ս6�@a^����l(�l�Ѫ�ۮ�/�2��d
'@Y�2����[mYC�f�4�Y.�X��Aw�����A�E��\��@��d�+K�m���Y����A�F+�6��~ڶ�8+֎L�)��{*�����;3�Em6��ߖ�ѕ���M�8.b��W�&]䦺���~��"����*틯;nN�l�0���ߤ���|���z�Q����r���i��0��.vˈ��:^Q�d�罯@g�y�ӋM�jѱ� K����L����?�Rb�;���G1Fcw��n�
8�Jr7�&oӘ[������S���<B|�<�wr��\;���]!�Ӫ�ܪ?����r�ҍK��O
q���f@�����ڱ�(��O(��[���ȃ��<>Q#�X�8��Ta�l>po���Uf�"��*ݦ�L�=�S=z�/����mt	ޟƷ'B� "	aY�9�	�٪���F���.�=��T�J�õμ�AFG�ħ	����2��`����i��,�?N;p�H(fz�V�]��kL����<��5��H���'"ެ�?��e�h��yl�4��*���7O/S���D�l�%q�g0��)`N!T�6{H7Ma7�nJP���l��I����<(>Cz	^3��`#�d�ڽ�7��d��� ��;�p�5>�����${�g��imhP��JQ��n��F�TY9���TWJ|1����E��\��ώ.�����5�.���ٷ�
�zޛ�T}�����1�P�[���d���: G�!^,M�<�-���ĭ�s{��m>'��OH�����ri�б�0T	+=r� �bҞ��0�X��L�C���O��9{�6��Y?�~D��P�vo��j�1�GΖ���5�S��D6(��/&G$�2�Ê�F�O�*���<��rf+����-Aj!=��Q
*<�����Çd�[�+�z�y�/���rJf���Z����V��/� �HERD+�7M��%��$`�˺5akP�^넁#Z|�K�$]���� `ay�n~5
i�ub&���_:?�e�����Nv�]���*r g���p���k�/˨��`~Z~��������Ǫ �P�,_(��+�Z��g�'���^9�-36/��xu|��q�oh��d��(x�u71���A�!�>�k*!ΙŴkX��۾-5�)k�E�k�&��鋠%[S��C�,)݉�Z��V�ݻl�<�W~�ŵ�s���q��aw��h�k�XY8��C�!9���
`akz]��pb,H��Y
/v�;(;��X⨿�ye���H��/�i�ɧ��P������,'<�bV6����ݺ���z�=���r��}���0�ob���k�j&���������-(���L�l#PV�����g*�;���"ɶk��q��܉}<S��Ĥ�l��]����1�S
(���Z���L��K����)��A�ζ�U+�O��<5�G}�j�l}�Wu�=�������y⦭�)����<�^���C^?*�$l'���,�����K@�Q�m��=P�.�df�W���48��7 em�o#^�J���>��1r���g��p�h�"9����?~4��ayj`��~1͸����X5��͋P}��A��g:�%֝[y�G���D���s����V��� �\�#��2��0ծ���TD���Xh��be������d\�UYD�5�x��W_�x�g����b������ 	F�RD󠝺�$a��viO�Aj�\���hQ 2>U�bdנE�dk�>�%�w�N�4��-��.��Zݴz`�O`��ӂZZ���<�$�_e}��b&(3tv����O� �-X���������ny3g�wE��u[��ڽ�W>�@`�{���d���}�C�J�W�Е����f�gq���f�E^zA���.ǌ����qq햢��W�����񬍖�%�x�3{�8홡���㭓g����S�r�1����E��}�ʷs�ػ�2DE���H����3ԇ;3��D���r��ԑ�g������$��)끡,���چb����ć�MZ�I_����A�� ���zFJ��p�#�癐���`@��X�bI��V����g����j]�/S�{���_"!B�����.@k٠��m��rKw꓉=�VF9�]Z��O98��߲���һ��!��Źӆ�FùZ�a��N���l,����-=��㷀[^���L�SQ����*"7x�|�֧���e�����@̳��Q����F�]�'a�ʃ-ECz }���t\�R>��R���2#�c�$�{�(�P~�!���xNV��`բ�[Y�\/���\���>���n|���[����#��6j3���'�T>��r�V�� ���֯����E��p�MNi͵�~���#e$�t<:,�.��C�}Q��;��j��5��9C�Y��!E��n��G�Vl��Ze�nW����q����wF�M�K��Y�9|̆�����٭�B�Zb��|�c5at��]0�3�D�ĸ=�w���M�W E1�{�:����3�z.�Hmp����x���cɳ3��a}�D�yQF��_�]� g�v�^��uy:�����O��K��Zw���(��o�i��E*�!y5��vJf�R�#��j�8g�����0U�ea�i��:P5	�O��X���%chR](ޮ�d�#JI}��2���B�n@�{�� ���Y+�J7�g�AK��M��!S^�ƨ�Z��")k������m��Ѵ����勥�q��XKV�m�G �ӗ�&��
�l-b&��\b�2�����7f��HzZ�P�^VK-u&�]d6t��d�\*����H�!�("��*��`�߬���P����.�I,	��HƅR�I$�UM:����!v���W�f ���ǘ˵ ��}�R � ۶�Q�b6�y�:��L�@۶G�Vj�	��J�E ��'�X�-S����~y@���0��Xe��D(ev�4j����t���p7��3K�����=��G4�4����u|?�į����.�.�#�Z���=�>��LT�)����MN�W ����LD���6u�L�D=�6��S`��CVQ&������^|��@?t�U4�]��YRO��=;�D��-d���+��vy���a��r�o5��ɢ�&Ê����״"(����Y'��.�{�G���{�dW+�a֥��7�' ���\� W	?ًޓԵ�=^��_��OX$�/��l(�(��:���T{i��%f �5aiL����&�V�i��`AgԀc�]�� �)Y!�Y�N�?����NW+U	>ܕ��Ϭ
�!l���XAUf���3%\R��j��r�����^JW�ɱ5��M��VT� ����v13��Q
|�i�����WЖ-�W��B�Xv3�(ٳ�Y��U�U���:7���U䣽H���1�φ�q�b�.�m{�rQ�P=��p	L��~�R0�m@�K�̻x�/�؂�N+�PT�5����|Y�N��K�:7�_=���������*s:XN0��U�l�G$�^�;�NXK&�k���D˷���>�k$x��1�u#_��uMs�H�a�NHG�?��C�.��	��j=3O�GrY�>�1�ԃ ܝX�̯1��Z�qo'P��9��'��	ƍ�wIl�f���x��]7��<l�t,�����纖��r��Ftu�.�GD�l�K�������'`E���d,D�|b_���Y+�1���8@�~�N��_3C�`~�[�}�`I-�u��gD3����vS4ԕ�0�w�x�\�ٱ�8;�Li�ò�9+@x�h�����Kus�+�Po�m���B׷n6�E*y�_`��K�-t}Է�ޯ?E� �MP�%��<�w%��R�&6v,�d�'���d����b�Æ��~�/�`3�ۍ#�cg�0|:.��aN�ٕ��j#-縚s��k����S�d[=��"/�]
6����9��y��*��!���`�Og >@'ٺʮ�����b��9��f��L�4�[ڂ�#�cg�A*'ؠ}��n/�K�\��M6|�z�v�?�����E%��C�?�p]e@a�@�z]����.�! @���ƨZwt�S��:E�9ZL�XB�'5n�����Jy���Y�N<9Ԩ��Ƭqݻ.D�p�Р�@f���z>0����[[���F��ʆ�G5��R�D=uf'�3���͋U��A�ﮉ�Ά\����W	�$7��w�4 cI�*�����2ٶ��q�u�y,;h�m�N�]V��i�)�m���ra��q��=�V�d;��뀞.$3�<�|�K�P��@N�NH�huį�*����XX��\V���CI�r��s^p����\�Ai��F3����!~��:V h1����S}� ݹ	����I�#�� DT?H����XS?�wH�LM�������Ato��Q�M��i�LاmOM��.�=I^� DO���]�,5�3UK�4]T�rϣ� ��b���a�<��~�L%[~��)�� [s��b��%Y�Z� �2.�ۡl|P��j�JP~�R��l1�"�������ea^����C�;����擶�����s��r���4�XU�{�>�ݣ0o�	�SN+�z3k0Vy�F.ɾ�`N��P�J�n�:�c��!Ƙ���-$��$QN���2zF���BgȭO�S��&����'�=6�����J[&�/�<0��޷MsL[ѣ�ذ2�X��N�,��Mc��-th"���6[_��,*$b�k���������*�5�R0�0Kԓ�.�p��'J��Q�=��{��}� 9)�Z�%���e��ү��� �/������ù�7o"�P��%����P�:A�R ���Jx�����!�Bםx����S�q��3
��18'FR��.C�i��z6��PHh�X�<�����r���=�=��~OC57.��NԐ��p���k���>�l�w�n������,�ϜG @@����ơc*�ٕ����E,?����C7��b:/�1�@��Y��R�
`@��.�q��,���0Q�wm$�Y���d�r<S��(�B��� �lgi�S��r�=�p����fu\�%�`�yx?����'\��X�'4�o�k������&'<څ��8"�m��0Z�:��b������]� �L�m���[Hb��1H8�%XH�4�$!�1���H����p
�j���R�/F<���c���4S鰒Gxព?��S��8x��e�El��w�b�'k&�c���,���4.������B�H��&=�����tQ��H4�R~]N",��`6oT��.���M]/�Ĥ���SCx��tD6~�ve�+���Q�Y�
���Ռ��B�4mӗ� ��EX~��j�3�?�e �wf��72mYU��c1�˷	�X�]@[�CS�g����l����UH�q�J��)�<�(�w���T�׷5J�>�
�����Y�$ԝ<OK�"f{p\ԭw$T�Ygw�T��pX��U��c��i]fY��VE(+VF}���������(f�*ў�qNZ�^��r�4��,��K���¦C�Ӈ�� ��=�63֊�����p�.g�(f���j��H�q���w0�e�"S�yB:�{\&ג�?
;�6�IV�B �Uǳ}j\�._���T�� �=�wt^Y�fY�^�z����_��ɭ���C�7=�cd����q��9������;+�p4�ֈ�㝤���Sj{j3�,Z%���E7\�K�3�@�!�g@7��;����� �܌�]���en�7y�*;mړS��'l�$�3��ra^�[Is�h��'emOt�o�I^,��g:̲��r�uXӽ���%
���V�wy�.`�whHt��ۉ��G��4����@�?V@T��q�����&��RF���O��EUK�b��~^2�'f;�w\.M����Tےw轴O�Wzž��~pw!�K�08ۨ,X)�������}��|aS*��q��Y�3�]!���G���ׂ}֎E����s�0R��O���2!�'���)���xl��Q��ff1��I+�����Ru�Y ��!M<�Oak2�w$�_��̠w�͸�����YH�'3�*��4"�=���|�u����hJ��{��㫉E��h*�TO)`�P&����2���Se7���ބ�Ĕ|�,����l�M����H��6:a8nW�F�D��&�&�<�A��h� �K��h+��]#���1a����
ͩ^��F���=�俌���A�%�8��������z��P.6�>���(���i�U@h��B�ZߐؓIb٩��e'���
A�*��뽜��&'q�����.�N��6����}��VLbjo~'[���}�ĥ4���樽�G�|6�$A5n	���H!y�pq.{㇢bo;D\S���l��Qإ��B ��
[0�7֛��m���+�7�`�#!+��o&��=�Xgt`fBm>.j��+Ȝ��k�9�RS�Åx��sʕoP������^S[����ׂ���;|o�j�@'#�#���=3k%^����
����ER����!�^Jr�ܡ���p�q@��[�� Y���dD~�I�jV[>���6[���Kֽ�g����CSh�D"��2�E�yg�p�5D���%#5�U�t�N�1�䊷0
GA�fd�����唜�a�����X/++t��W}030���4˶��i��JZ#�G�¦ʉ�7�g�+��JԬ��������P�Ӿ@ބ%��1ۥn�b#��;�.������T���[	����B-�ih���GT�>��ĬxS��ĜT�ܒ4��5�7�[��Gg'*C���4Gm��tS��G/uv�t�E�P�j<�v�0�405��{~�:Z�N}xa
iZE0(�F�V���J`$;�ըx���'ܙe����4쁰��7��1uo�5�a�Ɵ^/�!M���'3�=Q�x�[Q~(�2Qq/}�HL�bR�j.��/U�3�;I��B4���M�6L%LD���|�,W6�l�w�ۮ|_X�[!�y��N
�<��`��Uu�^�ԏ��g�:���N��Ef
�߬ �X���$ym`�!�}s�T�Ì^y�`@�X1r��qf~p2��Ôv��@��jL#�r��@(���:�i+'@��+��^:��l=Ic���g{��a9�l�+�2�p��L��t����F��:4�V��pQؾ��[�2�;�ۢ:��b�ܩg0�tdZ�ec�o�J��|I����{���$�,�R�1;C�ߺ�[4�}Y�q+oB�y�^t��u�ߙsp��ISz�Z)��A\�"D�.p3]n�x+'_7d� �����H
L�T�EC�+�_'��i��W()#6� ��Xw��oe���ÌNO���W��G�÷���V"�Z�_u���z���OY�œE�i�/% aq�Pԝ�LH�������{5�Y�H��B�W��v�t�̤���VҀ��;2�n��m���|%r�)��/��I�� �aל���CP.�M�O�W�M��jX5�1�F�>��U���M��&:mPo�wTN��DG�:�,d���̺��(a0��o^o�<�ǜ-e�z�tf<��0'�9�K{��F�1| y�t�1�.����H$��IFR6��P�75#x�-;� �0�$����41�M�h�����HK��K&���ٖ9o7�n��|Sʽ��;z[&FtLf�'|��wr뮭�C�Ԗth'���r��_N/'�q�ቆX�2��}�W�s����MxV�G�n18X�&�y�����^�������Ĳߔ
f6�S���x���A�09x�%o%c�� W�v�~���Uw��|����q4i@�|���;{!fN�O\G�r�O����8�ly�����bw�&���mT���b�ǡ�#���^R_9�H[�Аݪ�x��H����Y�W���D�,7��t�$�)���fb�s���P�y;����'��"Os�#C��G�����F����{�����j9,�x�Ż5,�������}�lJ�,K|�4�7D��G��N�h[��D/k���!?�yˇ�k�o�JI����L ��Bf
��Q���L���k�ax��4�U�5x	�?�ݭ��x#Dy�Tߐ̰�T皶=2�؈Xs:%��S�lJ����IoD	�i&������G'[��j�O�ds��w��dw��eK���G������3�CSFE��s+ϝ��7����p����&��glU""Ws�tC�߂���mx��d�����l��)^�J�lm�'�u��aDϹ7AZ�����P����?�7a��j�=<������쐵6��	�N_�>���W��	�"fm
�3D�SV���N�n����U&�;�����<[��Z�45|�a˩����}�z�O�(�$8�ܫK��k/�����r�CP_ �gAZp<K�k�
�<�	��j�ߡ��:f��t�f�
��v��﯃-XQ�{������ٖ���V����?�%A��e��#�7ޯt���~�鞮��CH�L�N��0�Ә40]���	HA�Hj����v)�V�T�fS�z���}��!F��v~�x"����̆W6�\�7_bG�6C"�heY>k�J��uާ��,��@	���<��t�׽V\�@��t���m�;yFY���"��~`
��<�2�*��}���Hvl�1�=�[b��y��m��}Aٮ]�c��ƯI|���A��n�������ռG��:����-4�Vg�"���%�ᬁ`�ipJK�⾡�����/����͋�x~�Yr�2��]�g*a}t\�+�_��
�������J�m�L�����G����m�lN�l�� d�Ud݌���q�-'Ype
l"��	ۥ�)}]���]Mr�U��0�7º���)�:ƻ�e�c��AA�T���\�&���'`�v��'�:d��H��}E�^0n�n���X�� i� 5���å��cؔ#QI�<%ß��Y;O6�ޟZ�'�gU6���jA��������m���%��j+ٗ�馉ɕ`,���r��f�K'noZ{dS!�f�����2�u�7Y����gbe���E��ٯ��Q�'�l�n�M5y�k�T�+�nܔ5�gZ�� 2=s�c9�у�����kaz��i:�Wܒ�?�l�F���NEVq��L���57�~�ɉw�Ǘ�"�*���9�mܣH�Hޥjb�-p�<�M�E�[�e�Y�M��=���Z�e�*I�Kۭ�?�6���L�� m�cm�&��ή�1�_.�T�����!�fɜd�s-�DB�	� d0��vQj�k4�jt��!܎<��Z��bS��_�`�~@G����^�l�|Ѭ�A�%A���J�a�Ѷ�!�|��1K�~2�We��:�d<t��5?�''Pա@`�y(���d���;1K[���'f������%�@Z��' <���v�͠o�}r۹1�Cݢ�pq^.��=�}�'1B�)4�p�P�!����O�g��/M=VX�?�5�:���aa�����K��ʹN����Z�uُ*�-y�����t���J��<�{�#5��%�����C	w�w �X�a+2>�F,����[[�z�#V}v	{�e��3�G^���_���mS���ȍ7��(�k��~�}
R�ӡ��s!��֨'%�x�������m	���v�Ï�z��0MK�E�j�_/����5a辟������ꨈ��3�Bz�sȀ�x�/�`c���.;�P/3��RM;-��1�+q��(�,9���j��<�]��5O��A�����8�ڬ$!�ѻ���
��P5�����E��f���\��9�q�4���W=��#$i�n�U_'�K�S~XքM�|	�E�h�x ;>��;*�s6�o��ݨ��� =(�|��ϛ�#�)$�N���StC��}��Ԍ��M��c�[��_�U�͓�Rݛ7�w&��5�F�l~Q�t'�x��]<�Z�wȘ��i���� v��t�89J?jĐv�aGXdsQ:Z�v�L0�]���C���_�Z">!�5���G]
k�L�Ć��; n�bLu��ױY�UY���#V�h�a�1gӀY�@v�Sr�#�k����ԗ`�Jۖ�h+�,�Y������b��?]�:�e�^�ȧ٭;
XW����="�Ld���i<��b�;�	YB�^���ہx�qYoA���d�S_8%�ȧ|���!�� q�E�J�ǐwQ�#�,��z�/��E��f�z*E��po�B��g���ZPN��c|tj�qz{�Q�)A�|��9�����Dx�jRI�ʚ�6^���h�lKU���L��V^�z�:(#����d�q���7B���^`�M.u�wN����]M��+���+_��;0�sR��\���z��}̻y�N�����7�u���l%�/�g���2ߡ��d�4��j�+J6A}>\8/:0�v`�� �*���/bo���}��ge��l��H�ϕ�y�D*�o9*Y�؛0LՁ1��J����}�A[�G���z˛,����r`�>a	�� du�������|^	�?�����]�T��F%x�/-N���]���EYv����P~�s��z���J�)��S� �����*��^���[b�:r�_&8�����3s�_h9�fk�X%;yu����u9c(qꡦ"p6c{��I�O���n(?[�<D�E�=��j��ީ`�9q�V·x�h��Û�G.�R�s�Nc6��C�%��	�x�1X�ps�	�p�ޕ�`���-V�k��'�EQN@�����Y��Ԫv�q��V�0W-��5ֵ�������Bw8Ä�.dތ������#8=�����V���Y�� ��Y�a����cZ�t=�g�I��E�-�^6
�c~��ݺE$�ث���yow߿�.�d���(g�pU� ��8]^צ�:�.�t��`�.;��d;U;F�s07�ch�달������^S�[�v9(A���t�l �j�sG�
������U�m�oh�$W��/iu��i��!�P��ؚ(3zdy���i�Z��9��ɜ�n��뉨aL����k� �xi��=M�����-�"!BB�����*$
c�T�J�ܢ�JhA� .�kcf�4i��:��D�4F��������W�v�q�����aV�cν��s�ku�n?½��%1���4���"S�o,Bú�D�zP�)�}Z��n��g������LI0�#�#]��pg  �G�c���Z�|?b�#�$��r����io$����^�~^]�� cnѶ~j�9pCTٟ��4��z�J�?�����}zz�F4T�i��ic|@o�Y�
R�V8X��k���b��Bp��m��ͨ���eb|�����j y��æv���X���_�F�XAw�WH�t� �%,K-� )�{�8�]��4oŨJ[���n=h�X�Zn_���G�2���a&�w¨�������%?WU��&dQL
���׎�������Rڎ�)����tYī�^`-P�C\��F`;/2�x�F�'����Nx_���z	��� zq�t�#�oyMDu��ZL��~R���o�N��y:��������N���,N����!�k�c��z�����bplR�
�W�DH�@�`_)�Y�@����U ;0�r����VPmX�r&N�ݏy�6*��a��\y��Q���� �kMu���
D��H�u(�Z�G�E<��gs{�L�������S�V��#�#�,�m�̄땯�ٙ�/��e%5�RXÐ3�G�� ��Y	�=��`�,��3��%�SL����E�{�u-D����1` ��;37�;�­+3��G�5>���P�>1�"(�e[����~X3Q�T�q�h_��wc.�#%�޺����p��5nQ�2�0:������o�Ma���y^��[��ϣ��S�{\0�� _8,v��1�yP�B����"�M'��\�@�4&�K�b|� �G-}���|�qz0��!Juee��џyMܑ���+z=�^��	��{�V���V��U�&��2*찏��e�9F���z��9��C���﹢͗S~�Ce�8�TK�v������ե�&�-��F�P%꽵��mja�Y��c�5��� ~���nP0C�L��(Qm��q�)1q"���ň Z�1����=�6�v�z���h[��Bג\������[�M���C��L�ֽ����/�gX����-�v�Կ�'�l?�3��w�Q�ŏ�@)�R~T�`�9����*Ɂ�~sV��5򳮐��JE2p��䒭����c��b��I�)��R�Lp&��v�|]5��g
FsXP%̮�����u���A�^��.%�,9�� ���)�&�Aح�c�}D\�c�o+�e2��e7��lݰ��	1%��9Ĉ���A��p�0._�I'�t�sc�B�v~���kac��?+��z��E>X��k�nTX��vEdL�a)�w�%��Ģ��<�ų��3
	�튇�8(ކ�j�r_���]���P�H^���B|��8�=bMt�I��T���}���h^� Au򔡩�g�]"���=<��#���$����Զ�������H�I\t7���0�,w2��=���ۣ~��q�T�=o�93��0��d���E�!��>�S�It��ň���䍁��Z(��������`����f&��?�ڄ�����"W��{9ǘ�W�6��OUu>�XE@�)��C`G�n��1<� �������xa�ǡ@�r�ʃQ'@��R�j2����򛠢�{�?qR���������ґ��JR]�n����. �G֢���&v��������?1�]��â-�
�~30vޚ�u��qG�ge��evb���,^��٨G�f =��U0��m/�c���fd�FX�g)_NKHG�@��맸���F~����j����'؉�W�^�8�����]�P�UV���=����M��`�Qy��$�Y|W�u�|�$z����0��GD�^	�v�1oN[e �C'�8�ި2=�jwN>,��񛨼	u��m`|��9^ F�Ϫ�نo��o�9��j�<�2��`� 垚T���bH7���E�$n'�~y�߄�s7�{�.��U9��c���.K�1p� �������wQ�����jGl�h��*�L`c�6Ԧ�8��v��5��=�l����\��$��D�d���Y��V;zCw�9֫��4���l��҃��_ʝ�v���H��A�{(�Qtr� �cL�Hۓ|2+�͠_�"P�7r͗��h����3(q!�ܱK�4��I��st)� 桛�">��'L)>��������m����g�}_3�)�E�E��7A�,-Īҡ���/Ì)��8ڃ1����ۅg�9���f5��������i��F�VB	���<$�ɀ%�M�%���vb�Ӏ��ǣ�~�%��/ܙ�Z�Q�[a)g��jƎ�^��Â���_��}�G��n��n�C^6:��z[��αA�j:l�q��\�0�5������7��Z�G�������,xg����u�}	98�t#��򑷝�*p�p�Iڼg~���l�`���"8x�������zm��'t��twV�������p1���[w,��D�^���\��AY�%\FģƜ����z�Y�朼!�&�]���R�q+�VH̋-u�����k�	Rb��u�jxh���
�!$�Q�:�	j�A��=En}�RL;~B 47f��+�71��mj��T����I:e��xȔ8@�S�p�|���/
)���U����%)��~!�������?���@�!�U�ZȂ�Gy|�\i������T�;Y7?n3�Qs�N<WR#{�Zl|�v��S�yZ�d8K鷡�Ob#���;f��p��o���}����-�=�� ���M���ʎrF\��n���u�������h�!,z
A���^��V��w�N���}.��j&R.y"�ϗ1�Yʵ�'|ѓ`j��Q�k�����W%8����<��p�B��t$�X
\��o^��bH��[�G�zw�z{`��]ƞ.�R��=���[�xX2L&>�@}WR�}�^}�\��'@�1�����p��-#�h�㜺�2�c{!'��Y�I�>��'���k�|¸c��r��v4�j�O�6l��du̦L�@M%"������@��8rhx����q��!*#YY���i޾�}�=�̱`F�f��B��~!�r�����dW)�[	��[�����R�1tT�P���y�Jl�@	��^�ܣ�j�� �+KxAx���Ϙ���c��
�L_��	G��3�k1I�bA���������N=|w2��~v��ޔ�I�>%�I�x8���9x��p����DU�Md�����9<�4q�h�Ku��XB��D*�P{�L�`�u�n��	�K���D�W߷NHסW�7�)�hء���&49*�4�/Tp�}?�jM>!�L�Dr�tm�'-\"��u�yeh�I�*--�K
#�B�(��c�.z��%�fG��G�b���[��@ ��\DkB�=�7�t��|�����5M����L�~^���E�5���$����1�C҂��N��q������z��o"٪��6.G��"r�<MW�s��X���$�D�E�wE���t�&���@��ALr��`<�6�L�W�ܱ��#=��A�V2�0N���D�6yd	���*�J���`���a����Z��,i9�W���'���;CJCFA� 
v����8�g
�e�^��o�����&J�!�("J*��_������	�闰v�y �II�5yۊ��j#j�~�.(!�V@�w$�2�[5:�/g�����1�F�G��e���Y�ҕ�ס���D��S�T��㫷k��.�`Kꋰ
%�:�U�kr���ߊ�~�f���yj�F2P�>���H5�Fg2O��|.Ws�SUEkp��˓FA�Y�'�,%�^ s�H�_�
�_��7-6�s�>�e�SWE,���!��H:�cפ���Z��Unv����;�Z�H��4�q+��3u��*�<x�d��=�3�f��r���-z�u� ���G�>��x)%.	�Mc�HW���ˣ��Co����Ցbu�l�>�I��4\}�&( �p�\����o��i��秾b٢�"�5Q7�����ˇ��Pgt�7ɞ���f{�����$��Zj�4��S����u��I"��h"�j��e�I��y���'O�`���3ԧ$e�ph�C/�5�eBd����ϧ��{G*�3�?���&�c�-V�(�>��aR>=�ȣD��*a���֥�w�P���e)].�����s:+�XM�O�Xul��j��2#�?f�qe��7��vK+�vRH�; C�F�ǯ@lLa�k�¨�!���S�L2?����ý��)�Ո�LH�W�7�� �F��\��o��kA�|����	�X�������l�pH��?z,Nܚ�/kf	���J"�A�u�� 
>$:��ٹA��=zĈQ	� p�@���O���FG�W�����x�e��v��Hg[�|2�h5�낀<A'��i����Q�w���%�I9ym.�	1��pݴ\���(G8��ݛK���S<<%.�G�RW]���ohØ�^��7۳#���QOSNyƠ��e�ƛ�I�LH����ԭzAa�C���K&�ic��!���%����0ї���wV�&E����L�;����X ���n���]癗�]�r�Vn�˩a�JՊ$<{�[_�0?��D��������^��Z��:i�Wz��w&_�S��5
��9oA?�����$�u�9^i��q��X� 0B�ia�JQ}�<�^�IR�P�ϓՁE�F�nIp6b��o�#�����M�Ň ��"�9�uв�`z��� 4C/)&B|¹CM5���Nz����#��;ƀxQo2U�B�;��5��Dl�����,�(j�Z���%Gq�kqd?�l�����%>sS�(`�b��VA1����&�
G,`���
4K�݈"#;�S��ER�E�{�З8@/J^�nq��쩐2o�s����m<ӛXLn
�&9[?�r���%xw>�?�	��2R=� ��f�e=��w��I�����ϦCD�l�R����(Y3ɯ�<%�=�`��o[+�a9
������vS��r�0�'�^�q� ��GT���..s�[ѹKI�L��]��=�!XR��<~�j(&T��ܥ����Ӱ�:W�^��Vi�70ҖN���3b�$o�5h��IV7c;�l�>�Hbq�6{mZ�i���y�������yV	�D�r��T��Y��H�����#�9?�S�)M�n�ɿ����##��}���9��'���1���_��cj>�������MD�P��sw����spFVޘ��^�H���;���"��0y����y�#��k�(��T��@�Z��͹Cb�AHք������`
�	��A��Y1?A.�D��eF<�N4�$��«ZL"����q����/��FHA�#�@�Gl��e����k�j���E[hv��nkj�$k�Z�EZ{��9ꉮ/�s)��Q�$5�J�Wn���H��3/�`��F�N؁>l�1��若*�A@Cen�~�dpFh|7��/�L�f 嬦lC)���{BT^]��\��3��-�%�ҍ�r���Z��e�L�;.Ȗ�n{� d�V�TG5C����<93H�Ƞ��<)'�����ǜ����FC�u_�Õy8>���4�|�`��1��n��弪��9�dy��#8☢��F���Y
�j����=4@�=V��HΝ�v~N�bO`�@���dRr�����X�"8=a�YԂH:��:.��\��p᧪Al�شj���~�!��s����C����e�ˠE���X�`&����^�����	������ⅵk4e�H:x��.xJ���k�i`AU^�&��
փ�m����g8`2H�p���_0�`����L
���rCs5�ޤ��:y	n��ᇋ2��( 7��z��f&��ʺ��̣'+��P(E�q�ݺ[�aX<d��~;\t�]n���|T�̙86�׊]�6�l����hk�)U��Ft�z�l<�n�;>�f�i�x;Z�/����s+g�{�������j�h:��@�2;�n�
�d���ޏI����G�[&��/�7UiHe�![s���}�k�Y���E���;�$��q���ȝ�:h(e"2�F`w����uQ�ڈ��;����i���ߢ��VRT�Fcf��� �����]a� �r�%d�P���X�@D�_Rq;~�O���[�<�
yk�L~�v.�����%����\]n׀�tqQ�Z���E�!3#�9V�>{0��Z	t�t�n�:f�Nxm`C�o�J(iZh���������c� ��5�+�xHPn`�TJ�1��p�m��Ys��#�sVZ��_����r�?���5�+p��jM'9�]�mP��(���=(A� �\��$�.9�K���� |�&��׍�o��]r4.Y���(y��<6���Y��+�c<�h�Q�C����M���#X�A���H��^�_�F�����(�na���������������+D4,g'[MDY�c��|5be�J)�}m7�%o�����[h���%�_Cȩ��9U6c�Ő��S��7�3H��$���M�>�B�zo��1G�-Q>aG��c\�4C{�!U b���%��\P}ǭ���Q�;��x�;�8	ů�0��6jT��7��K�8ԚƯ�^m�,��8��T+�����e���[v���a�ȦavbR��Y݄��ǳ����)X}�^f$*Ft38�(�J�AF~3��!��d����ߊ��I&��j@��"6�<݆�V%	{|�dJ���x㰣=�5�~��Z&dT�L@ue0�#���<r#pլ�đ�Ű�U�9���Yv��8 ri�1V.6��N9~�,��;[u��ڟ?�|7{�J�1J��W��n��a}
Y�Z*���b�5�`��]��>��<򓈅z%��A�� $ߛ�n� �;��nd��m[��Z_a6t�I��E���ɴR�_la��@�[J��v�X�����]�u3N*����$E������K�ƂJ������Q�:��L���K����EM�t�a[���lQ�8��/y����:`��P�h X.�f	e�Fs��~���-�f�H��.���י��d�L�����k�r��������]��.@j֮��ݔq�3��4Xm�a��/~u�]���$\�xH+;�
=o�,q<WŔ6:�v�չ��$��o��Z�	�����2۞���z��s�
�����ɶ"8�E�I���,�gک�����*���e�m?#ʕ��  ����̦�*p&�E��I16`9�ò�Oݻ�U��i����Ǟ���ܯ�զ`Q9&s��eS �r���p6?%�I�a}�Y�u`�0�F��>WH�h	�N�h9�Hq����k�P��d���*!���C�H"�24��V=7�[�`�1k2��^n���������Q�>�||�z�mD�;)���n*�3]�c�q�ԝ��{[��!�X"�?��	��ZQ�hO���,jl�(ͭ[޶Xh#�g��N��oi���޶���()&�X5�,�/͹����~�܊�餏��u"c2�`��T�̺?w�C|X� ���;��0%9H_�3����MB�&���f."�{>V���	�`��,�c��~Tز��"�z\p�K�Ѱ�q���ϐ�mc�6,u��u����zС�H&�!�G��PE�OH|�y� ���� �	���N�Z<���C���i�����[������!�n��e�H4~�B�j])/������i��45�z"a6A�}w���O�쾵}E�g�����
V���*�O���lV��j��6�xV�4�iKn��63�dm�"w� �R��oܸxj�� �����%��"��'G��<�n�ve�Kl�]"�ݡMc�)�(�1��A��_�Ia�}G2��m1����y�#�ޯϭG���1g�ӱ4k��,Ӕ�d�����p�F. �Y�h�kM��(�EO^�N��~�����"�}S�ǥY�dPs�g�k�Q\����`�_R.5�~�Y��)���e݅n�/���9��k��`��g�|�u�����Y �!�(z�O�8}f�����(ٲw��0�|-G�e|��aN�r
 nvU*�W��x˱���j�� :3C�� ���g����@��?�l7����z��w�~�ą-�}L��Wn�	��c���<��V��8U�B.�#ܕ�Ғ$�W-���,*"Fk^�3��<ш0��FhzV�b��o*�
��4�����ZFY�)�����ɂ�����;a��U�	�@0�ju
Q��I�٫�"G?��y'��u���4a�,� n]��טK%`�,��-a�f��]�[�*����qٲ5����+MC�`a�gf� ��Q��l��e�S
���շ#eG���u��+�ـ�\2;k*!(C�~�r|	��4H��}k#澷�K���f���Q䐟>p�v2����QP��iْq���u(z` ��B<�X�����V fjVh�݅�k1��@�j��xMM��D�/>os�0<k7��,Ѥ��k;�⌕��潪�V횀�[I�i�Zq]:���e�kĨ�낎����8�M]�w����f����U{u�)Y[p�,�!l��!�{� (�g˚�N�ZS�p�XSg�Y�|Q��'h`xM��K�<[��?fD:����b�� 2A_3a�nt;lSd}�3G����>'�J+
��G_�g�e�r~��ͺ��Ys�Lң��+�69|+����;�;�>\_aє�:��4�� G��D%����v�c�z�ܛy�[ ���4�G�͝�#�"�|��9e���w�f:Y*n�����x�"�s1�;�=�!��sZ��6~���5m'>��}{Ao\���c�!�$+��n'�w1��{d�u|*]R
	~���%�6��p�#	,�hf_�!�y��vK$0L���
�y���L'H#P�;�g$;�"9�Q�nOИ��-���TwVlbq?H��|>D�}"ri���3����Q�U �ZX�Uv���SE^{5�E$�{{HY['��x�c����3�5�~W��N�-��k�/o"�4�"r� �����bѪ=U㤜�� �+��eA[-�Fׇ�>��#��7j�Q�c���Z꥿A>[��]|�a/1w�M����u����h����F��W��u���=>1�|Q����^U{���1U\ĳ�H:��A�T�N�=w#9�Z�Y/f�O�|�����w'
;��T�7�(��v0̷o�m��gJ3��Fv�K�@��!+�@xAm�;��������[4`��Le�8�:�l�"1������̫NB�T��Y�s�Ô�@�?\l��>�o�A�u������.4<���GWi����Fy-f�h�
�ZB0���.�����,���=p�m���{^�%6��j��&�{�!�Xxg�{�
�1�:�}�W�AU������������[xP��P�N9��$�\�U+���TQ����.��Y dœ�t��+�r��\�aP�h�p�g\��m�GWi2��;|�ĕ��M'lܥ�Jː���'��7-���]� �9_O)	���ډ���e䢓ItG�ط,_�=��7m�}g
��ʧUL�����O� �`d#Dw���X����[/����X�PI�	Ͽ-��
��V�@�`�⿇:��Fo�K_��.��TK��!�:J����7,Ц��3b��Ƞ�	��}yv{^u0�`�#�H��a�Z�<,�1�
�xb�~&�wi�C ���{rϱ��`~�L��-Q-�(g9��кd��ʔ1k_ԥR��1>6jQ*a��etw�4�\N;���NU�]���ȁ� ��D�q�O���+rcвx|�30���͡%YdG�R�5�Q��ؼx}*�B�F$`Q��_�W3�2��MH����;Y~���.*�O3͛i���f`��i����l�<�w�x�� �P�mY��t̔uj�Z�/횐�,+�28x�J���b4pYȴ��Y������e'oc�4���6潗�p}A��c�2[���?�Z�=�1���k�������K���9�
WdP��п�9�.����F�Pg��꺤�P��*X�̈O�9��9۾�*+Ɛ�x��5bQ5re&`�U��y��Lt�\�79�ܫ`/��o�~��;���C�\WO���YP�Ѭ��ks%*��s�sq��`�`s�(��<\|���1E�"���Q��Կ�PﳣV�h((>��@K޿��7��(�����8��l��@�tf�(9�N¨:�xJ���x|X����2�q��~M�?��H�78�r%w�&�JNt}n�5⛌�%�)v����� �)���gI����aʠ[p�cM|�/��@Y"7��h�nit�̟����ؑL	D��A@�w�Ѩ�)��e�#�u��{?�>�\&�28K�op*�A���w�Oh�Օq�$ct�a ��*�nO���\{�uj7�]��=�)�+*�w.��5yj>��1.��b��z̊D�#���{x���C�R�V��^��\
���yaL�oز7�=�xr�Y����<�)1�����Ik���8Kk��#6���B
d�bo�1�wY�z/5���J5v�z�2y�g_�����IڝXnN��)/Ɛ���'n��"`���y�I�]�JL^������u�.��˒�NIk���K��,([��n�`������+I�I&P�󿜬M_�=���l�g�וn��y	U���Hԟ��MHZRo���|Ox^(x���U�F���6l�6h�=h�n�U�c���h7�]J^��ZcGa�#0;�t�n���`V�L8flQ�U<�H1d6�Oي:���K��P�;�~ч�K;����]R��O+��n�wsd�A��:�b�D��F�6�7���wlIں��/�Wp�X��tә����R�V��c��P�e�i_�1A/4����9��U �3J���`�jƦ�Rc;L���m ���c����ش\2�8���]��A��r_�'򝁭��F�~h%G�V;���hi*ӏ�'WT/K]��4�b½���Uz��$�����������Þ�0�b�ʷu�	��0�A����ՍNc�I��K2��sp�0>-�`�	"n�|���Y�_gt$�{��tT�讜ȱ�OeXA��F���Z�%%����a�7��C��7�9���^n���n��o�ԏU�r6g��!�o��
��!�OȰ#�B�?�w��E�?�HD����[R��D�p�Ǫ�ÛM����PU=^�3��]��t�PiS�'ڟ�b���L�'�`G�|L�GFcp7
ٲ7�۾�H�f𪢈Y����N]@�h��E��v��ZZ~����"�Ba�	��5h��X�L��#��`�8ڦ��$ɫQ��S�d{O��z5<�������_��R~;��ӟ��c�h�<��jm��\�٫Aĺ�Bt��62��%�T�ZQ���p��+�s�q=�i/G&���~	*���[{[[�K��`�`Ŷ;%����6�ʵ�� ]�kW�m�3�s;��A�3�q���Q��,�7[I��%k*^���"�Ϗ@�N�&�����!�����o�3 ��R2��S/��ӈ�^I���}�`�˿�����u��;j��˿,�L= ���}{���@�g@�"��{�a�y���C|z�yO�� ���[�'ܝVݍ6��r��%� ozC�p�a�Y#�H}���|����?H[�p;�B+�ݯM\�j�7�C���ƅ_��q�fy�I��߼�O8��!���+���B5ϴ/�<�G�{�ne�b:_:��������i���<ĲQ)hY�K��o�����M��aL�Ή-�T���+��nc�Ew����XS _z��k��������*�n^�J^8� r;U����;y�'`�X#����n��ໍ��x�b��h�\|9t����m���SD�Op��ә�Lf��ؐ���X�HDc���쵮:{T
:�$���S@>
,^Y&��;>����iO��G�?j��G����+��=n������;&c�3j�ן�Т�vAr)Vg&��Hƕ���z*�LI�5R�`,G*�� �Ľ�#�Q2�7�{�Eb�t����G�׽���"��Q���ė���>mk���	�V�~ɣy�B+���$�UR�iyU��
D�-�ŧ;���z�ީy�����T&�$�'+>M�?��hk�v����@Rk�+�Ҷ���t��9������}�׼,�ao���j}wU'�����[0�*a��2��T��qʛ�>Fa�Y穫��=��93���Hx��h����ۄ�yx�,g���`�S�	�T�01�5!H�%O��+8mO\���|������δ�ȕ�+�v�,����0�"#\�tV��\�S�h[�w�"����
L������*i�hӖ��4��u�� �l����Z{׍6��c�� }��׹4nu�U����C"�;������#t�	J�§�l���:��m������\*�Aȿ�P՘�J�F�G7���/�C��y5�v��6���/�E��p�Vy�xn�wi�L��;��5��)��J0����gs&v�n�Q���LP��͇���_.uu�H� a�]�!�B4�h!��Q�;ۿ� h~>�\�DPALz	^ڢ3����,�_X�NPɥZ����}� ��Hk�Y�G!�,I�3Y?Y�T�] �����c�� ]<��jk��E���(�AT����$�#j�60�GڿW>�v�м�S#�{NDS�T�04���k������5�j�@�4�U�b�zQRV5��	����N�$dz|��L�p��ܥ��_*}IN��Z6V9U}�hD�-q� �I�ܡ�=Da�{��U�tL82h8(��B���*1L6��4�KX\�S�R��fr�&6ٮƩ���gFیo�^ﶷ���з�f�n{V	���¾�GD9��X�H��TcD�	�-nǧ�
�w������V\=��>�ԇܦ���\!+5�o�C���:F��i���n�����y�<�@t�����48��W���AV�"��K �hߛ�c�v�H�`D�������A_b= ���~+&��]�������ճg����� cE}�� h Xgt���*�Yi��>@]FJ��
��?j�s9����d��[�/�Y��i^Dֶ��{����1#"ҩQ-Oh�C��k������������'ԏ�v��׼H-���rQ9��f������h���.�W��؀��[�>@]bԔ�DU��sI�T��C�L1|�����������,%���k��F��yq��ۙ֦�^Z܂f�A�$Fd�;�o���l���\<�4�+я��
U+�ǚK|	r��޲�Og��eno+�h� �,Ӟ[�
���pp: ˧\�I<n���8s	#���}ן�o}��,�����������U����-��7)�;A��������b�i�b@[����i3>MQ����Ɨ�(�
�� vxOf<�T ��Đ��K�I���R_q�`�7�CL#0�OT_x�f[>fX��8����~t�	�P�0Q=^Z��i7rz�
�Iݲ�m0.��gb��DtJȕ�:`j��Վ4A��m�V�V�7qf%/���*ѡ�=�LSޔ�聊�k����1�K�-�r�`y<.�1m��fݬ&R��(,u��+��U��S��e����,����Q��)�Uł�_D�+��"|���";Ak�'���,a�"�8��K��/��W5)3'Uy	����|r���{
q4�*�u�R**~A��F��6��q?����3����['���G�)Z]m�=�2������I\���d����f�P��M�'\�2�F�\��(�gN�� ��P���۰��������z�qS�}��<�B%���d!���G<ДԹ�0A7�\y9������������f;�Z6Av�;"c%+��ݟ��m`F���R§�[h����/�:�i��̿�=As6τ�g>'�{3Ԕ$�l�3�<�<����~�*++H7�ƙ�x�J�a�Ǆ^��p�R߾x�de��>��5�_�/%-E��2���U HJ�l7���~vdT�;��I�ʱ�O"#v>O����k��Z�s�_H��t�
�(7���c�,FSI'7��U/�2�x l�_o-gK�P]��b����t�du��o�B��!�h2[�٥���Z[�����g�D�R2��c��@b_ߤh�@|W����c�V�#V�]>�ɑ�ޖ�C�t5�Tk=w�fmu��!9QOL�Q�^��m��r< v�@��Ec��~�%:fZL�S�ܫC�n7������du��J�Vkɵ�)*��	#�J�g��79;j2K&�dV-Qp�^�Jm����>�N��6/.o/�l���	�%(����"���=i�;U����#�}=V"BxQQ�,;^S���� �Q[n�+�����gA�VM~��d�#�s��9OF�?�vz���]8�r�鹒FR����c�NT{�ĕ�_��ǻ�T��tU�?-�!��sFRX�ۃ�0�eu����c����ޒ�XC��k�3����}�*[/��6�4��n_٣��Vo��T��l�U�o�ݓ���7��֕��]�l�ń�rLܓ���Z��e�&�S�?���K#��%���+K�7T����,��Ք�b(�#�� v�Eְ!z?\O�� �48��˦b(~|Z�����b���}�]��q?~f�Bm�rR�Dɺ�I�pJ6�鴞�q.q��\�3䃷�N�e��kJ�c��i�A��5�w"6�/�2Ԝ�Z�8o�?2�j�
�
ؤ�%o��6l�w����A��o��lhJ>�NrV�i�����8���A��P�;�D�;������:И��S��z��dZT�Q��
�5�˃)����,q�$|��w�5��\���WGBR�S݄)�<����༯�60���Йz����,��kEx3��G_4��'bѪqw0On��T�Ar�����Рz����%�������!�^�}��; 7T��x<�����7�\��IANY|搒�O�7M3LP�p�u��Aӕ�rb�����:ʊr���OM��,��PG8,�]3�a<��2Rخ����(3o�VN�����SA�:��r��u�� C���E7��M/y���� �(��x<�Q�l��1��[c�N2g�i�q������0>���hZ;ȵ��Xu�]�^�E"^�Xy�@��y;]L�mO��Ԃ�nt���/&���A�숨�2�h�8A��/��ғG:�C#�3�-��q�W����"�.L��p�O-���E盃�w]�7��mQ�
�)���P�HY����@���4G�wv����L��J	�غ?p�c�M�,i�#<�ą��B����MOm
��-�ti�0/P���5���_� �y�MM	�`q*-�i�����g�Z6,鿅f|.��"�ٷJ
	<�����	�6����sYi}	l����̅��AHg}��*5ZR������̴�`��\^�%��ڋڕ��7�!���6�9� ��Ab&B����S��g�;ȦK�����P�A��:>g�"�WZ�?\σ�r6�ۑđ�6zk�
�y8�3_��`Kgʈ��=ؑ����L�z����W61�^C�U=��A�7AǗ_R{{$î<�ީ��d��pcOM[���w�i�DZꀶЂւ{=�W�W7�������!��aq?��&H�k��D�,$t��<��Δc���]��oU�T�� 2}����+������a5[%ttG=�LT��l6;�Ͳiz^�$����W
TPf~!�q�+}Н����V��Q��E(:�� ��oT&f4Cesˁ�� ��TC�T�+ˠ��{�Ɉ)��V�b����'�G�N����tT����0P>nܲU��ѱ��_��Ɲ�{�����uY�ϊ?��wT5�&�g�J��=�>��"�#[�8�e�2�F��@�2g��o�� ]R�g'�ǵ�y?[�#;u*ћ"%���*֜Ķdޏ�'�p/gE�E���^Je��@|0���v�/M��H/�_^�h�����z;��\�9��l"C#��3���?H �pys�r\0�A?�v��(;��}L��r������o��b�D�_7��)Ι�4O"T�֣�'�I����yأw�.q+���(�P����r��!G�L��c���R������'�/�Ƅ�S�ن��\��A?O��IJg����VZ�̦�|$�KW��iz��L�]�0��/X�b3!�,�,M�)`Y�Sꣷ5 �85�͚���>$YpӍ=Wl,��!�y���7e��fT��-�G�lZ���@�Ubz@������������*ҝR�﯒� 4>O�Pkk�d������}ppV��%MD��z�v�%g'2�˷q��=Fi��6�rKD�#!�pp��CX�K�i�>{��Ld `�U.o�t�sZ@���C����X&��&�K��;�����Z���(�mA24 ��Dz�e��4=l�u�{1m2v�mI�Sr��ҝ�vC���{S�bW&�ZYPٗ��J�8Q�=ޮ�2��ԁc�ԭ���I��O�/x��-0r0ɸ-e���|���J.ІF������G�P]K�� Qdi�y\���y�D�s{p��[�"QP��D�w�b���0�����j��ДQòh�U��,P���r� -听�?1�#���T��X��@��Ǹ�c�ɄTYT�	�6�z�'uuO����R}Cd����������}��_i���-�{���1����k�x��k�Cy�#L=	e�������	���]���ڼ�G��~�Q�}��Y2z~Z�G�x-�M�]����?�Rɨ��l#0̖>��nr�z�5��g������U�/�b���K�f�l���1��v�z���m��L�>/̡Ҁd4���4M��@mr<�9�1�QZas RGh)
S��ú�gn\J\;D�1��9T���!�r�B�Ӹ
�i�FԆUU�i�`0����f��9��s�
8v���7���� V��r�^ȉ��g��ou(��:[�/$�u���&�D)�I�*8���"|c���'etn��{D��K�G|;u�5Y]�^�UR�yV!��v�'9X� (�,Q�%�Cq���G��!]}����}�yZ���+}u�����lOR�ݫ����m��rĲU����!|}��`�>[d�X�<�QRw-D��@Տ�fD�E�H���'�	�k>�3�/�dtW���ٚ���$�1���cM#�N鄘~�n��$�oK�/Qx��Vn��'���B�_<Y�+GJ�[���e�Mp:�6�K}��.nTkYX�<�����.e��p~,p\�ш�1T�{�Z�2{J��=�����R[���Ic*�*׫j���	l������ts�屚��ߓ$��4�x��F��̪������/�w~�U�݈�aC����mA^:�&�q�W�����#��'�:��<1�B-$�b:ͦ�\d,Gw#r�ܔ,;���x�g��6�m":�n=�-�6;J� @�=aVъ�;V6w�������3!'��� ���}�cm&�NM���5� A9�ֹ�F��Y� ��%:g�������8����r�|a��騁ђO"���}a�7�6�S�ܬ����_wd	L���m�b��Q�VZf�d�5\��8g�<��<2�=ݯ�mF� �%$E����R?(BLI�g�}����,�Y0Y֞F�}ġ ��``�c�.����"�Ǎ�w�G�FC �C �d�F>�E=�)¬m��$����)�H ��:$O���:VIo��E
�@��x%F6�;���ZI�	�Hk�"�?��0���-�����C���M�n	�@KP6h�h��U���o����(�����_��z��@L�^5uѽο�A���8kI��F�`����]I�Ʒa�Q�K�%�5��R���yd�K��&����!5�g���)�%���
����k���nd��_�GYr=S�X��3+j��~<���P�I>FOV2Y��V�Rd�v:w����yL��dH$#\Ll$eFP5@�����;���Z��sա�?�w��S�y@Dxߊ�@L��#��ߜ�O���a�ȟao�m��B79������Di�3�Sv�l�ز�ua�����0�8�(楌�vI�/7��Hx��N3�g�$�c{��'t�{�<K�-�	�|¤�8g����
�w����Hh��Z:�Jv
�H�V�Ds��yN���_@ll���0�U�2�E��n��VǺ�,գ�I��� �gh�\{��n�Z]�+vb��E#�J^�	�Gd�x�?&�7a=�al�#Vn�M�UV5`_�6!`s����t�����^w��b��|-j�㢶ͷ�����!�� ��	t�b� @�x���n t��$ ��n���0��b�zeq\�IC��q�w3���p���~*F��\y����mt�_�ʂ��iL���Y\t�[E ������ݴ�?20)���φO����𖄆����\v���=93��;)�'>횷�9k_������Lm����ȏ����\#����DZ��+Y��6!��\eŽLz֡�wД�6G�K�[^1|�2xgN�kI�Ǧ�X��Cg�:W'��1�FC}�T>�,�]�\�l�O�V�N.�i���Ț�͛���\=�O�$�}-����������R�_[�D����VP�:&ǏK����]� �i��m/�7(��=�ѿ��.� t�Ŋi4AD���\�[��생k�F��D@�
�싡:�85E��7�{��Bg�%���y}����doq������2_��7ˇn���@��Ww�_#,e��H=Z\F=���,�f<��P�af}4M��2,��u�>��b��?�J�Wcu�����O/c�E%.�}�/�����D��{,��_S�̢o�.�5x>̨o���>r�Y$�] �V4NWլ�j��:\gU#ܗ������J5/ٌp �����X+EKN ��l[Դ�ϩ��c�)�/��a""�4>��K@|r#�#�`|N��?�"�7�%�!p�c��)��9W��C�G.�i���98}��v���t���W�e ie܈:"9�Q��f];��w]�L��p��X����`�@;��'&�6l
��=	����ձ�fk��f��ME�|C G�^����H14������$+{��w��a�s���Uj\��3�B��+�w�K!��|�v��ۨ�5��vXj};!�D�QtWԳ�D|��,��^�D� �&�vB�e}xL̒�(�,�׶��"��`ks�1q��}T��I���KK�W�ڤ:����rh�X`>�6� n������\��ϡD����=b�t�*�#��'��C��I8��R���`t��/|$�3����%����~�q~��i)W1`+��Q�z�WSᙗ��B�*xS�@p�\"8���AW�+O�n���3�%uc�Ƽ|s0<D+�_O�x1E�r*ջE7�v�����w��r�˝,98��+%j�n,I�
WN.`�b��߳ �yG��t5ZH��ب�٥��$�o+�-��^o ґJ�'�����p�[ߎ]�7����6�~ꤊv�E�+7�YB�_0�ls5��� mME���ܸh��1rj��~�З��/�$-��q7�k��Y�C�)���>IջL�s`�.^��46y+�Ws䮁��)Жǘ���,��2�Cgh���K�2t?��tr`�(3���Ķ6V�H��c�!��p��߇2J��Z�p����3c���s�|�5h����Ws�)� Eξ��k�px�R�C��`�!�	�`�܏Y�������*�G��躀*��i��{싶W��ܘ�W������C�R�zm��/�������q(�Kf(y�@�\���ؤ��s���Om%Ę������Am��|��:��K]���ƘWi���U�ٷ�!;�	i�5�
�fk|��2g"��Z�u)0.���=-[���j��*�����D�.�Mf��L\i_�;d���1�YK�R@��1�,������%+ښ��wL�j=]D%,I�s`c��BJ����d9{��)���J_�K���'̯$t��qz����oh���ǟAj՞�Q+�)z��P���g�zF&�60��{��v�fr�m�~��?���fs��!������ ��%>/�{���C;I*;��H��ZW�Ƥs������d�,1?],�ۘ�$�+(�L�X��~�9J ����`$OT�خ����s%�U�I�FE�##A} �~��K��&99E���3T��ܻ��κ�_�i�;@��?�jt�i�� A+��#�,��*ᷚ�~���DE�7���p)P��E��B�m�'y���R�5�|W��`�&I���hW;Cm�f	;;���a��(I�T���qr/T�*>�<�v�1�.�r��O���?�v�+��o�����zΙ�pl$Ț��ny�t0�^��=��!O}�kTS�¶�_9*Vnn��*�8�$� �?���a��l}K%\�������,~��"g��ebw��9旝0Ɂ����~���N��J�u�v����:�{6sT��SҔ�b��"�׀pb�=��8��W�b$B4���c�2%���S��r晦�!n��4[�34�BV<�904q+�s���S-��@�"����:Y�D����ξy�>|H \�&�W ���k�,�fBB"{�2�MH	�
��3;���.�u����U����s���{Y��5�C>ņ(��7�y�����N�(�du\������*��畑<��PCKB��_葢(Av�/c�&�[z��g ��L';$R8�=(��'`�e�C���k$�4�_�^���N��Y��l��S�]b�[=�X����R9-���;�h�_�s�^��d(j~4����
b�i3a���<3P��j��Ô~*�u�Y��񯡪\���k�3���A�G����tg_M�Y}{�7|�n]ji����1-�Xd>��Ȅ�(�}(Mi�[5Iܝ����&��5�&��@@-S5L5�(��1���ZVYRLT^���sf�L(%�-ՎA���{.�I�z����KQc5?>j��pp/����~$C'�rX�|s̻��� ���SIQ�6�r�Y'�-<�q	�-{^�Z����jr�
\�"N@���"Hؤ�o�e��B-j�4vW0�b�E':4���`ED�rz�K���q?����ġ��3��2KH>��\y�ճ9���2�[]���!��/_%�5e���*V2!{�"ie�1�P��j����{���$��N�(3(�J�O�b[�9 I�>G��]��Z�r�|r����AUC�R��|�M�ڵܦ����{s�FB_:��|���b�$�Җz���Ω��n�k5<hᯐMM�oJgY�n�����%��� ^��Iy�{J�ٽ�"`�B��>����YS�W#4�fV~|wz%�r�e�� �-���X�ؘ�O�$K�� ���3<~��R���K^�@�q���,nA�Hሯ90njj�?�I&^1K�@D�"B��e%���y��
KI�eDg��OCS[����v  =�V��z����<�cE���+�)6ar ��k9�2�\N�ᮄ�j^S����>�]�^7��g�
>�4�D�u�H灘�:~����`G��K3����C��N��ڿ�!<�e����~ƾ�)��q*�����f�?jTD7+H^��E��X>	�cO�^oo��^i{<N۪t��z��~*���5ɠ�	���Hش{����l��(B��"G&S*�FѲ�˒y�0�X`+��3������G�������6���#�R|wɖt4�����2�鰽В<4�2�{1нt�D��Ď��5�'/,50�Lt��8�ꋝ��.�z[��r({�A�_���$�Y��K�����٤J�vP5�.���a�A�]�?1	��k
e�J��Y@>�*{�'�$����Ǎ���X+,�l�ۣq�g���S4�1"���o/���y3���K3�c����]mq�����SY}*�Ue�"?��dp�+�L�c�����@�G�1�kHٔ�����W>м���hDnM�t�-��R�D�r�B��0{�YӀ�mCF����-s�[Lj�zUq9>�L�%��;Q*��]9�p�̔赺zF�}���$�D �Z�(9��D�����po�����75	�	�e�dR��i}�Ul���_ ��/����;�φB"`�@8�Lz�
���Ŧҁͤo%�UH�&5Y�\ �92�NK`��T ���S�t�p������5�	�\a7�)�ú�%f�A\pQ������{�U��.�Aie���ո	�f���-���Cq9��lC*J�I���m�wו�]=��S~J���q�}	_==���I��"2?qK|,}&�I���r�|�ՎapX�|��sC82�t}	��||��db �7��.�G:hF�CAcdb}l5v�?aƱ����9h��{@��}N���K:��3�7CW ���]R)�R��������z���|O���5k�*�+�Z�χS~(�+�Z2x����[�/:�k�`��
��#�n�I���ǳ�'<N�j��� �8	pW�Gc-ϳe�ZV�������P�����&�:�3T�P�DC\4�S-~~��&v7~ۼ��M�+JX2A�W��t��ۥ��`2̕����[	��f���b}ա��b�.m��A�?
Ci��l��Æ��@�#.e�;x�$Z���#i��ڪ!N!;�utN��Y̔Ѿ�y�Z���.9A4��z��z�ɹxE҂���*���M��$=0K��< ٟ$j	 �g���(�nh�+�>�EZf�ua����e�I�N;@,��F��2���?\[ll�����3E��T�M�o�3���;�{Fj�R��d���9�&і�E �^��`��CX�F��m�3���j�]�7�kd0L��x�#��8~Cn�m��(wm�8�_|VH��.^�	4`�kN�ץ�3�Wh�v��UìG���W؜�=L�U�G"�	͌78�@���(6��0��*�X ��8���G8U�2�ȡ.�G��c� )ײ+�/�)M�?���{6�@:�p�&�jT�����KO���H$Zo��w(#�lX������~?�6,��|�=���S����#4&�҇�H���h�?KF>f�|�P����Mt(�6�3���xj�2�Ed��$eR��S����<����Sk�Yt����I����J��Z���5p�R�j�>��"{���<*�p'Q��J�fV���
lZ��O��-�uzx��b5k�����$/��b�K,�&"�*��g����2Ċ�H��j
03+��HD1:u#�Z�HaI��16aUE�F㼽��ՀG�e�� 4k[��Υ��굯�֮�ۺ	�S�\s���$����,��f����m%����	 �x)�V�Ȍ+#�3���<s��S�������B���U��wX='`d{��,�|e�z:����l��6��ѝ�S
����;yg���#ᲘŘNj5��(hf}�ȫؿx�s|N��Q�~�>�l��62�D\�"�9jɑ�J1�ܓ}���h�^[.����B_Y�
ˇ��$Xi��n�2�����z}i�h���@1�*�OX���!��ЇN�ރ�8��àPY�{��-MM�]B�˥<�n>�탈��RbYŬx�S1'Bg6Ԕ�db�c�S��J���7���+��q������i�$^;:�D��٦L�W�Srw�������<�cB'A�>�}d�)���y�4Q���{������ӵSG�ӧ��,�*)�]�Ч�������uī\_"�ee��M���Q��o%�(����¤XLE����>ʺm��hĴ�[��ۗEϑ����65��N��<�U��;*�g�3F�v�ɑ���Ȟ3-c!x���.޵�d���0���Wu���U�0������R�~U���N����=	=9�c���0p�.!��
U�#��|^����.���N�����gv�TJa����d�\��&�����a���UW*\��^�X�pu�C��=�/c��A	�>�'f�k��a�$�J�w-09�����]�{c	iG�J��@�?��`id6�b�����ʱo����ç�U?0����l�?o�R�:g���P��Zn�D�ڡ\���N<��.�y	�*��n�h��\����*�|>젍}
��iJ$���[�� ���΋�c4⒂&���AX�Tf�Ftd6
O�懮�z$:LX��Ǖ�o��Ȝ�f'�Ll��&cI�W9�k��W1�t��r�u�T!�`����f6�yʆ��?<�+$2�S��QO�����Ka3u�#M�nl*4��")w���5�W�c���e�h+_ YEP��`��E�����k������{������\*�� >��:��ߗ4��$5V9�s�T��U���*��d�\/�˗�F8v1s�!R�`ʼI�]�N�=ǢK1b�J�M����uX�� �ѡwG ���?�{���)^o��ӚUX�.���n�e���Ԥl�)	;h@�+p���(�q�J�GM�c�IT��e�����A��ǋ&���ͯ{xh>�G��'�o�j�v1��3ӷ)��zax�bRʘ64�����#����jh�<,4N3��.`q�:񦵕�2�*͂�c|�U&��ϛ2��P�2H[�e��M Ψ�
�ɰ2}��*���<�/�b�+���r��9�%g�k�+��K���R+�t�$%���&Z\#�ҕpt4S�'��\��K�KC�yC�W��2�ϥ����INE��?�Ez��a��OZZ^����3~:�-U��k�L����!L%f�h�t�f�#��`�H�svE5�8Q�D:2K��ũ]6�e�	
=�؈]S{2ȅ	�~}��{�'T�'ZG��T���fX����2��:�B������b1�<q(?	=F�j�_^;�7�IZ�κ���x0v��2GL��K_��g�w|p�������H(��.��ߴ/��N�����J{y|�"���5��O���BZ�G�D~�l���t�"UH�\�I6{�X㵗Â=��n��mᎼ��[��Xihb���$���C���@���9���e&���O�Ҋ?�:A�������&����}N4�j��|�;����~@9�'��C��U�G�@�9��M7i0�b�l��[͘Gm��a����$J�c��U�_�H���   �媄�t��BQ���0�&0dRC�J�n?��L+ɲ����H��@'�x�']�!� %�nB������КX_XF1)����2ݝ������Q瑱�h��z*��Y���G>�q3���:�tc�@�6��C� �FWj�m$25>�ҏjYo�\,M{%>Zy��g�H�c,��nf�>,f6v�����!b
���S�b�ϒ�=����B��':��S�G^�g~:�Ϸ��	S��8��13OUtn�����F�\j��ॆ����yD^����jK�i��U�}���
g���k���%u�i��_ׯOP�i�8(g�����-9���lx���Vn`����3���$fU� ��[=�+����Pi�������}��Tw��=�Sl�Ǎ��K4��Q*�);�HjA�Z�%"]yd>���tDo��L�P�B�1�r-���MzN�6Uf�:Zu���3ތq �F!4�i��N�vV9;�ؾ6Wb�ĹC�W_~��0\l�4G�eW u7��u^Lc��c��B5����0�D$�܈�Go�����0�{��S�P4���%��*��s��+o��e>Mt"�n��G��Pk=�"�J�:��"�ޏRܽ���O0Yz�S�(~����w%�����l��r��y�2��9M�pA����_�e�I}>�Z,�D/6e�8�b��7[�G�- ���r��{v" d��}�j9nJ�H��U�g�̽��hi�m/�u=#~L∣XJTv�iC�3&�׬�Z!�<Y�ԩvy�����`V�K��c���e2?��x? %B���O��pr��2�0ۧA�[@@v � �� � n���t��a�N^�o�N�uZ0Я�,� 7�9�K��� ��)��������肧,�4�"#�v�8[>v)�A�/�^!��Q�R��ɱ�#?�?f���ְHW7�L��bb�5x�z�WU�u30�����\�|+_l����2X�j��X� ���!_�1��N�i��'N��k|���$!��r�<��94QM�E$�O������4�jYe����g|FtI������]��[�ɿ�Q�ۜP�!�� ��*Y�T��^1x�9�иzGMc5+�4]1�@�u���8�����zi�����me������5���>O�0��c4�L�����\�`x�b��x}A���?t���+F�ȷ����/DDE�{~J�R�$_�妤�6���$�Q`Us����1�7��E�F.I4+3n���C�vR�!�H]����]�� ��{%�9�f�"�z�	�;TU�u�Wޤ��Vu!��:��Q�\�D)�n-�W 	�����϶�ԡəM� ���!�|d��-̋[.|�'�>����8��R3��^W�/�QZߞ���\s"��N��<�r@�i"��t������t��d>�0�(���*���)��Cv/_� ���0���M�(b�U4�3h
Mc\�=���,��W���]����+��0�8�I�C�3��.lۦ�p��{�W��+/<X�
9��Xt7�%=S��86����Q)>4Ԩ��OV������h@ #+E��4�%����U�_���ط���!B��%���(� D�z�	&��	{������<��+�2��I{U�f�ţF���k}z��-��$P��z�Ii��T�aۗ��I%C>�LE�hB�G��Y�b����̣S�[���w!�P�J�uLz�X[8�J�K���)��a��*�wΞ��tuuR�	��[2��d�!4��i��N"�1MM�W�-!�y��8Bw���Ee�g�hi�%���������p��W��4Ҥ=�=��K(#�����U�hڔz�ׁy+���}�P�]�e8\�E�"TgA^�P���I�8B��I���76�+c���L����l)�l]�o��P�k�"l�d&J�'dV�\�>�d�c�Z�����p`�"v�\�4W�^���,�cq4r'w��f�g�^=�'�}.� �n��/ȃ�Yޠ�ƕ�(&�W[<(���P�N7�=v��~���U���J������C�����u�$v[e���$����ډ�X����T��=�pV�/���>��qΎ�Wp�3��=
�e���Īz7�X9���|{��s����cbj!{M����Сu�h4P+�^�V��;����R�������8|1v��bM|��?gF���>����|��
����'#J�p�Bs,�"~`q���R�V����h��|5ɀ�J:�~Í��Gu�E�eT������m숱��H�{��p��퇭�:+_�3���*�-�X�r)�����
���z���k��&$=����?��x�:��_O�5'�4]�/���� �װO`I�.�����x��L	q�r�� >hܧaPa���4�@O-��^�`�H@�d@�WvK/���9L̎K"�x��5�⦦}^&��������O�s��1hl��c�.f�ӏ|��� �a�'	�ƯE�
|�#%�}YT���� Ox�UԾ��*f�c����tH�y+(::��YG0�-(�
�2�q�
t���GT��eT��T�1f�o�����H$ȍE�>m~|�'��ꘑ�t�"�i�[�v(bp�:j�F�q�=k�錼E�ʇ���)��_�N�&���g`=�r:�@9�~���'�M���,bA���l`p��-oVLm�֛�c��
���P[�HOTJ>6~�A��v��f�=��A"�R�O��U���)��� [�=Ʌic�q.'�+ߦ
���#�+r�^�w��[*i���LT�����L���s}�tlunCء�n0(6��m�"p i�:ӈ��A��|�M��Y�����˅ �΍��G.��3+�V�!����֑�'�ð��kKĹ�\���c<�ZDZ5����x��A��f��� ����<c����']:�,q��#����n�������{l���#�M\��"&$E�]'��Z��(�HC�}P�o��ɷ�$��H#���sE�W �1	��9.�YyJ�3/2O~%�O��Y�*U�m�����޴쮵_�p�?�y�5j���v9̱P���d;$J�O�}��X�a��=j�R�ķ�o��fy)�Ħ��=�'!Y��k*�$�[l���7���O�>I�^����6q�U[�����/��-��#M�ka���5��
R�N�[_Vв�F�~aDMxtF6�|"C�鎑q¢���D{n��Hm�G�$�qd=�7<����d�c�we|�ɺ3�%(�b}�s|���ʠpu�;�������dw�+�$��x�6I��<x%dO�R�˕�-ڈ��S��{�^� ��n�����<Gݡ2��Ub)j��d�-Vp}J?� �$��g�L�f�0���bw��"���DDĎ���t�&�L�t�x��aɋ4.s�B髯*�����g����ӆ���6�K���
���L!��YI?[e�m�y��9�cۏ*7��,�y�tuP���$��5ݬ�ݻf��s��h��
��*i�I��p/�b���|�Tۻ��)no���~~|��+�ދ�B�M�G����W�_P`���(1�ʎ_�v����XiAU�)�h��,yf>԰�F��$����Hj��pC�lk�G�?Χ� ���]���YE��j���&��A��6���V8��b��E���@hΖ#�)���d�t��w6�-᭕� ;� �.@;��%���!�N"R��h�=�OiU���FY�"���P���t4��N�u�h��9 �4�^X\�K�C�F_��]��y�==`O�&N���I��h
c��-gC�X-��,C[9ړ]���qhT� �'M9���:8h�M���En_\7rDR��}{x��v���D�Z�7�5W#�l4�Q�	��x��A��߼#(tOЛã�CT)Ѭ���4��ItڤM��ь�h0ϡ��?׈C�p�2� �]�l�����V�.�M���#C�+����|�2b�ՒG���$1��,����A$Yw����vS�׽0˪h�TpN���i�=��D��0󶓺JU������6�5��ڦC̰aT��>���9	�y�f��i�*�[Z4�(��폝�*Ph|����`&$j���Jax_��m��~ɬ)��"��[=-�a�4Z��/���{\�!��_Z\�
�����)�/�hb�T�2�`i~:���n ���C���"xD�m�#4 �g3�mR����ݗ&V�~WiV����"�=�d�|dF��eKXn�W���-�z�sM1��94��|GXIO�?^&Mٚ+�}wd�GQ�Ȅ:	�Fg�R�+)N:2�3�H��n�u_�D���ȧ����%?fgN>>h�R���zY�HE�"��|�[.U�+
�\�u�,G*b�>m������!{y�VL��	 U<Ťh����B��pZ�'�$����E^%gDXV������JL�,���R�H�2͚Es�5�w����\(�$��|Tvx�0�|�V���ݩ��E��J��Y8*��a�ۛ��&�����(��Q%��f�t�����@m-׶�p>f�"���Ce�st�I�zm�9�ǽ��&0�gw$�J�����#����c:�Y����iUc��2�B�)&Q��j���2!i�W3�+8Y���*���&�^B�1���?����X'�ҙ�-/���]�A�[sD~�с~܂�m/5wg��{.̓t��Z�n��}������+[9���x$�@bkw��X�[���eeç�wH�s���)����k�?�w�D����#9Q�&*�gpUF�4��S�c���沵��K'�R��X�FUm��/���<�)�� ��������$3,-bIm8;�W}�c>X �B�.Ӣ��>1�'6z�R�!('A��k�G2��(���:?`~�h!J��!�y�u��q;A{��c,}�JQt��W�
N�Sc^z�T���i���W�#�H��]JH�M�х����?�wx�Q�����]q_���*������8X��M�{x����A:qZ�n�'߼t_��"搶_^�)�٬�]�a�0OҾ�:&@az���Bn�p��~.����[xE�(��8a�'N�J�z��FB���?ʕw�f�&��L���f�FӕUH�]`G���r�whG@�~���]̢��}�*��u=��P��.�w{_1�cƊz2Ě��Yt�F�3�sg�瓫ɰ��iI��1ܥ� �o�/FI�uL�}�8�D��?���4����H�d���X��o"��Ɛ��o�����=	%c���^�?�'��:	0�	iZ+��մ���5�A~�'Ē�y;Zcn��r���C��E�$\�~r��`c�\���UZ��J ��r���Et��UI^�����yZ�b���[/��h0O�yT=���QN P�J��:�՝�Xܰ����B�h��i����k��w &+e\�=g�v�\�F{S���l?��X�ʹ���@jQ�[�����q�K~)�XŐ4�B�6���N���MN�3|�H��p�'Q�rW}H	3�Dwƣ�b~,����s���(�a�]{,�a�7�,Q�\�-ZzH�o����qm�w����ZTSdΤ/ԶV�Q�C;\��U��w�T�@ r/����.��Q� x�jL���w[�`{� OZ)[�m ��E�6؉�t�A�"	�m��^mɻ�y��
[Nb�+]�T��g���7���4�ʫө���dP�AC�M��:9er�N��G�\�q�U<�0"��aW<}�Ppy0V�O��쮃X|w5�Z�'�H1�3�r��
hK��;�],����c�b�s�3�A�J��´�}ҷ7w,��<j���'u{E�s�+�u����q�߄��is����m	���#���]��y�N/V%���[����	c
�9�FX�ڋ�R��ѤN�^=W@9P� �k6e��+4�,��wE�&p�Uc�Tyo� �ȃ�]�}�j��7�M ��m�آ`z~I�E�|���b��GD����h��ֹ$S���� ������{�����r��tL+����]�^L��o��1{H#�u�PS�����n;17E�\� �T���QU����	�5��6�N� .�F�c�Q���b&�LV��!�*�?�C�"�^,z�9#T��!B%u��ښV��T����Α#m~�Bl�_�H��֐�n�Ǧ>�q���hN"Ir��bo!��n�?���v"��Q��O*h��B����F&��F0B���vu�NOu�O�sc�F���
,y�k#�?�a,�}ѫ���<����J`���9PdLTe�[����������ArȄj:7�<su�x-'W{���Ӵ��3���P�J
�b��1�A��%�}� ��T����n�Dt�EP#��(����,�X���iȨ�֠�~���9Q���B�������:�4�"wD�a��P��p,İ2�h:�c�����`\�B��Fv��c���.�~�J,_^ō��E�T�	ۺRV���z�����8��d��R���6x ���ެϬ��e�fUz�v�ĕ��W��( ��u=�:o��=�P�A�S��C�<Mh��=N�|���J�O~���1�N�H����gc�jd�~t�p��2�n�'V�����u�*��t(�+#�8KfQ��} % �ϡ�`�J���{�z6z�f@�2�#���eY��n��E{�q�W��D;Px�z[^6�4L���̯=��[f���W�?*5��P\�U/������Dn�O�.	�rs�������+���S|W�)@h���b���?[q��OH�v�I��QU|���R{ȡm�\w��KBx+i��Ri�A���S����_��g�wc늑"~>���A�J���Ҡ���w%�kd�
���Z���P���A�&�I�ԇK�'656Kw]Y��c,�qu�'�����4(6�n9Q�uP�CR�?��t51�-�fD��7/�u!y'�����x�k V"�7���Y@���gDg��Y���w�����1i�����8
U�[/�u
B���F2�5\��S�'��۪;�8������ZT��e��ib��T��d9����K�[�J!	�<��9��o�ҳ�-��bR���q�:%��Y-���aG�g	^��ln(ს[z���� ���+�T*v��.1�XM�p6ʠ��]��F�Y9= *E1e��]>&
�N�p�.vO�0��r03y�>��M���s8�PH匣t�#<�����l��:`q�� ��*k�#^�����	y�	{C�?��.eC?a�e���,p�qӊ¨���|�W�Z�x�w
�P��i�EMd�l>��L�[��hY���5�k���d��)�Y'T�JPU�tj�躝��Á4{�p�VD�nc���¶R�nw�X!>�l���l44~��P1���6f�|����vv��M�u��V�H�'����y8�r�srW5��~�y�G��- �׫ލ�2���̻V�-�V��A�tpB7iW�|��Z�)C+5`��'f Z0 2!�w�x3iy=�^&/�Q��/
�"l[��9G�ݿ�hT	nH�(�0l�:��9�����pK�uJ�k߻�Xh�6�=x]P@fH3gUe,�f�v<��m$TUl�g�m�.{X�#����eU�-8
(w{+����?3) ��w�З"+������YY(�in�-�?�x;�H��@�Pi�.����l������VK	�i�0��(�̅�a�R1+�2��"	�٩~����k��%[�4dd���v�J���\>�!?����iv2����C�Ý�2��
بsI�č<s0z��L~���3�?H�پ�K<(
o��2`�S;(��6=���~0Ŋ�]V�t�l1���0~�sú,�9�%xo�\�^�f;̃���~L�!�[X�X�0�\�T�jt 
�R�YdUQ~���T�n�?�ʻٸ�cEЗ��NK������R�b[��!�,�������b9�� �^A��T.BΜ���t�M�<
�*�p�K�	82 G��\���@�֜��;EO�[���Ɉ?�y��Z� �I�3���-g����4u�zk���X&G?��-X>W��cx-	"�-aDp#�OIVWt���٣N�\��o�:Zµ{mhEq\7��&p��"��&p?p��u�v����R8�gL�� ����UTN��kOA-Oƺ}\�ɾZ�m��)O$���#t<y��o|0���F
 �3�ոھx��6/�=k�#�mL��o:[_�x��Ȁ@s�c��U�����_���^Rn�����<����꜑)�7Ӿ7¬$�e����C��3M$~�G��������6������ �����2�����{�Vn�TC�D`�{�2l��@h��62v��)�UrM�Q>�0�o����x���1QǶ�V���߅��� 0jK׎d=N�� �L��k+�7|J�2���0����A���ݜ����^o:��Q�KC�5-A;`T�D�OѰ��V����\ulO'3���K�y�ʯ���,R\{��ա�<l74�r�2�Ӽ���N����=�B���Gg�l�)�!PBg����n],m~��F��B��2���������)$�ܼ�G����7w��Nݽ�Ö��,�[�p��]�'*�ħH{���;��v.�
�������jm˕�#�|�HM�_U5��V@�X$㏷�wRl�������kp�����ůcT� ��l8]br����F�.�}f���fYa�u6��R��zY6����C6E�+�i�L��Kg�73��2�6m���A�X Q�b*�C* -j~;|�$�-/*��(��H�&��
�,f�Z'�U<k�`�#��ញL��.�u��omP$T�|z�Lۻ
�GN���'c��c���2 :uez�ș	���k�6n�7�j�T��c)����gyy�\B־�@�7�v��=iVC�Y=n$|��^%a�_�u~2��b��Hl�����g�܌��l<R9G��	e4eW���G�܂/}��Z�f󰆖v�~��)/7Z����G Od�1��qF:��(�ב��N\�6��<�ߍ��g��'�0_UtC)�{���u�,���JᣳRx��R�����)ۘ�O?�L�j�,onE�4%]��b�~X5��O���տ��l��p)L.�
�KP���Z�������h�*�=M�v` �~����K�to��m���JXj��0���hp�$��� ��
�2���ƣ�ƑyѢs��r��]~E3~��1O@U�괾~1Mи���XՖO|3�8�8�j�8J�ŵ�V�G�E�m��2��dpz�9]�Z�v��Q��4	��+��.�Bkо*%�d%��7;��t��3�:�dV1D�������ܗ 1��b���'J\p���I|X1�Ù�L�N6Ll$��;Ô,o��P{�4lP�}!���eC�z����5%ݾt�<)�A9�8�Lpm4�	,e#��i��[�
��9��;v��֑��Dt�f�\ z�l�+��o�T�����%w���\=FzQ>���#����x�R�*p��[!#Z̜ì��J��s��8P_�_�l�T��E�Q������O���&�Yw�]3$����@>h�����+��� 3�SsEF�F^�Ja�5���VND�bDq�>�3E�y���e���r~b�yG��&^��Y`��#��usw�y��/mq�|m#Ͼk�-�]�`����3�ђ_����L� ���J3R��H�<��������8�u�T%T���>����*�����,+������F���c�o�<Ǯ��0��E���TM�"F؇����.�.��c�uɫ�m!��K"��3�}.�a|���lֆ�O��'D��vP5�h^#OxG�gq�������01O\tHr��#^I}�22�����p(C`�u
XI(g��ʧƳw��F�����?R��z�؈�8#�]���.�.�7/�n���2Gz��\��p�{[��t]��V��p���㔷畁��~aԹ�F'Ddu5�w�5x��s㦉S.��#u���EJ���װ��E2���w�^�;Ɛ�P�TF[3&x��e���N��$~+6�8��>
�?�e.e�).�AaA)M-��XXv� M�ہ.������!��ў��A��:�5����I�����ܚ0���1e�}�,�kw�b�
�z��A�Vb��isx̄0W��s	�b b�sD�w����8������24�5�Y6 �ͦ�
��� �~�p���XO�-�B>Lh�~L�mf��D����㡋M���>�p�s�(��]��@���j�T#0ځ�p��eU��,;��8������X�!�t(ASr���oGd����C�	����{�~�Zy�nC�2i�f��C㙘ā�# �1���nV�s��.�f���6t;|SX����򖪛$h>K{�P�"�er�v7�$߅�9*6��=���r��7\y&]�h{������\yY�dKq)4���.�������ٟ�'�i�]Y� �#�^�T��&4����AF���>��m�n�(Ŏ+�C�����m�V����JnKHn�;�e���)�V���@�H[�T��X���WI*���Ӹ��
�\�����^�}��'%f� JB�ӄ���D��)��E�\X�:Ƈ2+ׁ��.V�F����%����BcL*�I����� !wϵ��
w�N��ݏv.ёf��#
O��6����q)�'��?���b�����&�⩧�$�����b�5X��e�C���(�q�qS�� ���nt�|W �F͂dԾ٢��f�fk=ޞ~[|���ֆ���0��/��ɵ�D�����w��l�@�r�=�o���}���f�Cn���$V�	�Ew�=�Z��9l�mS �A����n��`I7���o�6U�n�7�ۂ,�Ly�V��7�g�6�bF{VD��ܱ��=�_r�Q��uUDD��͈ڈJ\�Z���r�w�W�Q4�3�`���
��)�(h`����s�b&ՙ�W�2�Q	9Y�1��y�"�R�%!�R��(,T�c�ku�}3�&hf����$=���&�|i��䲸'W�P��Sp���p�y
/��+�\�˜Ϝ�ߎ40�c3!Ur�n�S$
��\�u��L����QB�F*��%�t���]����8� ���RE�����i��W�a9>q�i����`S^��ƛ�F_/D�8~�p퐼3�*u���׬b����>bg�a+߆
�ك��k0w�@�Úٺ��!�L(h�sT�.�@䶴9.�شF.l���x�7�ી���m4�%���D�� !�%�B���ˌ~��h:aW_҃��f��+�\h�Ŵ�N����o�K���L��E�OՂ��6�A9A���@��i�M�[��~�8)�D��A�該�My�`L��5
,�ߥ�C;��=�H���ɫ��w�6m�*����o�XO�'R�V��=T����������m��K25z�����Sa,h�UC*�?�Ȕi@&5q�Ǐ���dP��ef�%��$f�_rq�w~�/�H���Ɖ��v�8���w.�N�3Ukl+Ls�4��`${lӨA��M��'��y��x���rp�q�')�P�{0��M�n����E�)�X�����V1DP�S�F1�	/�c��KeT�W^e��PŮ��d��M��⭎j�O'^FS݅�QJKG���LhrE��/��ୌeW�e�	5᳥ϵRXx���W(�e5P�cv.��:��T��&� x5�-�\|F.�2��U��Za�SK����l�#�Ͽq��2�:an�l��2�Ӿ�����I�rx5��i��2�9M�Ǹ�]kg�H�3�)j�Q[N�#�=�7��Q����)�B���~D�tͮ�W�SFޟm�S�C>ʬ{+�w泅�`�����L._��z�`PɒqX�#3 "�ʿ�==�F�4�0�!K4TE��^���ʳ0�Rs���>v2�`�/�����ye#��ryaON�j��T�����:c.���!_�w��W͹�ɟ���Do&T���%WX�N�;�&l����e
�b��8��'��iW��ڢ�/��k6��r���M�/�;���;��n��B���|�g۞�8�d�x����j�p��YƤ���c�g�ŀ^C�	.*�ػ�������魯���h�_Ep55��/�;-�$43x���ἐN$�ڠ�@^Sw�]�?�E��pf}y�V��+l���s�u����t=�A�J��1�q	��Q�����@$0+y�!�q�:�!�/�i��{"呖�_)๻�%�g"H�]]c{EDX��qϩ�>q�HO�bV���Q�ބ��e�c��%�P��<�I�yC�?ڇ��vkZJ�h��k��1L�%�;�}�zO��̨�>`�΂hIӸ��7Yb񝇞j"���?z�n��y=P��L<T�4�΁��G�����Ѻ�W�f	�Xy��~G&�/%�H�~ИV��0�o�[.s�=�_%�#�At[��b��G՘VKK����(6+�qO��8��n)�/��=(���r�nW�I�p�����8�mo��f���Q��4p��G��`��r�-�Gk�=�=Y��˩a(^�͇���;��u8G��D|
�\I|��Ʈ�v5a��eŸ! ��A^��B&nT��u�]��&����N��X���݃�S3��x�GA�"`�T��R[{|�E	��i�#�2�}�} آ��sۥ9�N��(߉:m�i�F�ߢO5B��Bm�)<{=z����2ڮ�Ծ�U~Z��!�y��[��P��T�t�˺�ݥb��~'!��3�+�oX�Oi�B8yO?Agtg=�|Az�ҁ�<K\S�l�^lC�Y�K=�Z3��3���LI�>�fK�2=�K��d<��w���Υ��q��ng^�w@�	�m��LSݘ���[�i"�ɷB��� >b@��p.��k�cv�k��ƶV���9 b��̜DCB�\��s$%�.e�_7s]F��q��h3<	��[K�w�m�=~k������f=H_�ɵ��(�bH0��@U9ƛX=�m�ygy���� �(�<�i��?}��7�aG��'WW{+��fW���	�*�_���~��Ɩ��{Wq���p�򤥅9��E�'K���4�Se�n������]�5�k/S��|J�
GF��S�pcU��4Ո��w��O�W��Sã-$-&(�C�������?_Zh�D��B�pya�=W /�PR�:� �>�����P�SqPS;/.fr �ml`�̂H�Bs�D��Y��۸4�m��9�d���N�C���Wq7g_�_����nx^�����vP��,˻ૺK
"�=uK{�S��W�QdA"��|B&��N�b��^E�rq�[-����|�a^�������(x�|�j��XkC�T#ʵ�y��䱗U|�NH^m�ik}|��M~��vL�6�z��v�D*����-znTQƦ���^�qa	Q��Tk���0�<]�~�	\�y\'2�?��%�﯃\�_v��)���]#Nh��� �va׷�k��b{p��D;������\K�l�N��n�K���7s&F��t����o������_W�6et[	���_g|�y���,�tT�L��_>����gq���(��,3#X�o�'�W���E �s/ Ǡj�քo�+�G�����
5C�]�hn�zec�,&ÉD�v�B�5E���6\xV''|Qb.�٬Q�ѝ>^�`~�%.p��IPӋ�S~��6�F��Sc��1|恙HN`�F�����X!]NԤ���O�� ?��3Ѽ���Gqtq���g�R���G<���Vt&<�-j�6�;B�{۶�b�h���s��;�9���	c>H��е���.9��	E9{�}��G����a��M�ʤ����rc�J~�FԄ�s�翻Gx4�J�\�-�ӵ!k]�F���%��,"��G���cJvg�I3�UUA�;��/B��&{ż�ǋ���apZɩ��"��Ⱥ���
L�N�Fھ��`J#'���~JX��N;�`%�*�� ң�R�����C��"\Uq
˚�f��Z̲��fI�ΥqmU���E`����n� �m$$�ޘ�Tk���!9�<9�j��=��_+Ǣ>4L�K�<5��h��-?��z��u��j�x��$ǝ�,ibIS��eݓv��-wӂ��QqiA�Bø"��C9�zBJuw���3��$���:*�����N��C@�k�.�L���#�W�F'�e����H*	�w�X�����O��A�^>N�"_��~��U�*5�p�<�[�JI��(Mf��F�	�.�����0{��Հ�d����uFHS<�NU%�M��]:1�-�V��Ǝ.�?ͬ��C���a�}-�~h�*�k�ɻ��'�����DGT����y]���i����d�<��/Q$���Ԯ�I�:�V#�-�+{���V�5��F��-�p*��8�ىJ���t�[�\"5���)ӟJ��Y���fi���<� �+��V����!�R��gD�J�.��+f�Ʒ�d��u��_)zA]�+�C_��ݯ���)��(A}u�����El�D.���B�`j/��S
m������l�b���Aj��Xw��ʦ@;������q�mSGk������GAV<��m<�k�+�������E�/�h-m��a��s?��fڊ W\���d3���n��\Efc����k���؂�2�㫾Y��y�(�a&j3!<"8_��X@�z�7q�B%��פ�IȳtO�+V�D�9R�A��(��6F�l9�ڷ.#���b�u�}�%7�RM�+�݌A�PL�%�!�u,���G=w7�(��#�Y=�Ӈ���"��-�� �A�a���!��;�P���EmV���r�S]�ip��~EP`@�I7�.:p�f�1��x�cUש o7}�n)ǈ��v,إi�e2�P���i�e@�xq���M�
����ގ�5{�׌��t�ݠ-�?���娞����T�9�Ћ���ڟd3w��ұ�;�L;}�F���*b��#��l��k�V��N��eN����*�L֙�h�|F�й'� H��}�m>������Y�Y?��"S�l�h����M{�n�И0U��}��-q[���,������8/�X�B�D�Rh�O��9� ���M�����l����C�&�Y�|7����J�x()������/��*%1GH�lt��Z	�o������V�^�l��d����bB�b@c7]# �(�����F��J��;���qBW^JM=���1��z�a[�d��>�˾�� c)��&)����-��8C5q@��ZPۏk��u�u�n��!-^�W�t���;?��x�9�O^�m�I0��m���K�3 �pՎFm��������<B�H:�˓ ��Rk��i�2S�/Y�]n��ud��N�4lf�Wɖ�%�5�i(=VY�
L>�|ӄ�X�M�! ��gW���Xb۞C?&����D�u�o|y��\Y3s�i�E��d�g��Y6`�Ȩ%��wMe�U}j<�?H��	>|yN�����3��"S>:�� ���V]�(k�A3ʔP�C-hd��_���Z�VL7��3SEo��R�jO2���7\�K+D1��~�%���~���[i=�1h8�6�	px�������,����pː?yw�;:nS��R��4S�V
ז�M�S�E�B$�7�L�4��f�1��B$:���B�=�A$�ZEc�"@����j�s4�rg����b�]�Gm�E�M��O8�ԃS|�������g�oA�C�jK�!��x����g�Tdo�ќ$]f��Z��Jw_���/�:ݐ���d�'�D
��V	{�BwƑf!��Z�#���|���3H�.D���$�@]}s�I��S$�����Y�o�M�Z�o2�`�/</9V���]��%�y\fH�3�8�������Z2!� ft�0�P����gS�]nkWp�`ljeH>s�ڲ������U�?3��߱���h�A{��냨�P��{i�W�.�w���fjͽ���S:��/iy�mZ����1����9�[o�բ������'$P����l��L~@[���|���[� C8P��J�Y#ِz���� =<�	R���ޖ*�?@�q���'���i�R�>������?3���C���z��9�^Ȯ/���+^3r�q6d�?^+	i�a�o</�!/`�c���chj�
��RyI:��>�N���"���/'1��I�9�y��ʲ��y���V�8N�����`o�3��mnۋ놫�0�]�� e��m=���A�ڏ<7I?^o�L�'X�k��(C�,%kX�+o>�V�U�N��\ϻ"<�7����a�ЖB�d�iླྀ��AA�Ck�
�
a�X3ꔈ�.�)�nę�g����i����+E�R>M�X,<[F�ާw)�ٛ7�Cm��E�0[����ߵ�dz������}%�~��b�2���>6�����-�B�2:�0�;���,z��5s��9��R蚟_wN]>��ҧ�e�=<��VRjH��sB���lg�y9l��D�;Jw������1��4Q�*<-�+wKƦW��^c)*�rI��|t>��BK��fr��l��B,�co([�6�eA�@�*�DҰ�𪜗���(<���<o-4n�U�y[�K�l���I2%��f^[�\h:t�h��j��K����@�����żМ\C�[	Ce� ]�=S�d,|2C�M����]�YG�N�<�C<q-��[�,�%��"����:�m� ��V��A��{T��+ҁ�n�����Bݻ��4����5�!5B��BE�?XX<õQvֹS��<���z���Ց�fg���e���$OG] 7���{Px�l�ӝ�Q���� G!k̚Zjh�79PG	�	���޽�&����s�N�0@a�(��E,�j8��)�m|8�	J����ٍҸ	�ơ���ל��iQ�P��h��1d�>�	a2��Em�k���4Q�w�a�3{,����=�<����*�'f,S�&(k437�(����{=��^��<�a��5����O��#s��w��娩R�WXwb%vj�*_GNU��f�7�$�U��sE�ƁT�f'X!�1��ˇii,G/}���td��DOil� ��p�0��/�O{1$���������!��kb��&���R��{ꁅ*���Q����u�M�~+�
���$��n���}v�(����?㲄�2z�Y�[��L���؍�!�V-r5���?!�j9�r�6< �-�#�Oڋ�v�z|�f<�A�|f�ڨ�%pg��Yݠ�y�yI�� N�(K�$�ߎ��P��˃���`�L��Qo/�7?��4M��ӵ>.�,3�_U$y�$'R�sG��x�R
9��Os4hQ�����Z�;�GA̝��a2;��c!���y09�N_C����!��!ހ�Tk�m�N����z�i�UU���
ïՔ�=�
�s�y�j�x��"��+�z&"��|��n h?+��ZT�)�zN5Y4���	8�r�-GXGc�u׺'1�E���hsA|�ݙ��D��S�e�%N�t]��`$�7Ԕ�q`w̭������tE��e/V���F��E�B;������W#�9��v���r�vҪ��cˤ�>}����vڅ���{ �}�`�i���i�O_u D�|��-���x���7��n�Y��JMܱ{r�Z����-�����Da�Jcu���4h�*���;�:������>��-?��S��b�j]���h�Y�^t-���]:X��a�c_s�ķ:hS�9sN�`��i���G�~�U%��v�o��̤Tt7��5j`�k+jY�]=ˋrI��2��)k2�=��ߊ��B���Ci4pn��� C=!��o
���M������KB��}���5I ��)"4!J�Ӹ�?ܒ/�Uh��.|ݵ�E��*O�Q��|�W��q6�LӢ9��հ�D�z&�wx������(ɛ�M1��
���l�d�E�Zo�j�a��@fӫ�5]$,{��@C�}�~E���yo4�<nbS�M�w����3�Wf�]�ϥ�QuH~]ؔ�0�_L�H:w���/��H���Δ"W�`DN�K[�>�(�g�����R%�O��	߽t,K��&��\Ę]59�Ǐ|�K ��Abe���~���UnFc�0����i~	_t�����ᙋ���辯�[���sty�����sÒST�\��)7��šH� �Y�퍱_-_R�A�dqr~7��������c����͡��>&,j`�mr����Y�jۏ
-�Ͻ�ւ���3a��_��B��T����JD�RB���m��]�]x�M�"e�w�6�4�:U��Vk�$X6��f�#�bȇpU�����;�����x��SP��.߆�"�s5�K_���̡%�`y
s����뿶��ŝD<&;8��f�4f�i�e��$�e�� >�D��ϞJ8SC������C%�O� l.Gt�q%�zQ1܃ܢ��O>�*y�ӥbX.W~SyԖ��{x�>�חM�n�iu!�[5��$�
{`$%mrC�[��շg˭��0�ͼ�$��ǹ����[e��e�.K��-$�p��
�Ep1�B�K�Qʃk�����i���N��)W��"�����K,���4\��E��M��d�)��-C���"��%0�Z�����v�܃|z�=�$ CD�(1a�5���+b�N�
��6r � (k����C��:��`�R�"凵9��IEpj6^�e���6�e?5� Q�1���`I�-��l��yH�C:j?M����ԝs7����Z���͟����K�'k*o��i��@�G� �jL�Ql��*�5!��������)=ݚ��q�<����8k(>x�W�Ol%oy�T)f�ڱ@�z��/��ю�rFHŦ}� �qE������^�ܾ�����Юg�<`f���D�]�ǳB�n9WJRV$��$/1\U����nw�<���~w�"Rmb��i�`0Z��z�+��
\S����M6��:�;�g�K����]�GΗ�����"d����o��=X/G�');��Ҹ�g��pr��b�.�\�~�c���d�O�O����x���"{-
���M������*�*�ǧ�S��a=����i��#��6��84�����+L�'�5��dC����}��0�sH��wsvw!ڶ<��p�¦��YX�n4�)20XY@��OZ�Y~�h�����;��R�,����3�I�J$u+.�߫��o���r��=���<�?��0�#����ڦ�B�$$�!�o�\u3���?ev�-`\��0�}QpГcպw�Y��0L��*S))�8��YK�R���?���rrҭ�Q�g*Uk�H@W7
�a�tXd���&W�r�j�T�G����S��ݿL�3M���n��� 16nF��_?Dܿ��w}]��W�i�4��\!����ab��;5f�/Z��@O<q�z��� �jFx�W���~�l/a�e�}[X�h�l��JW�/�jnB߼�j�oMi	o~Cb0l6B?����� �58�f��v9H_e�$�&{�w�?�xm��d��E{�@U���~���ԣ�VXw]=��X�t7�G�M\6��=ճ p�}���2X&�
�7��+�^�]��F���k�I�}L�yG�eN
�T�&]J�Y`*�oD�(܇7P.�6l��|>F�a{�FT�*?�B�]�gc��y4(0�H��e5�-G��7]/U�#�a@�ۡ��*r����Tj/�Ư�O;��*�7��4X6�|�z�2��#U�\��$��616��^�ahA����\T��>���YS_��-a�V�l;�b,7He����)b�I6,u�����>������X�q��U�h��B`"�5��մ��V\h$�EiH�!�N��;�i�#|;;"�}�ӻ�i�u�U�J-���8�� "G�斺k腍�����g������!���3��;w���V�/`{�j�4���A�w����=����656h(8�F�
3�1v���	��&�MX�����@b�'�E�+��?���@ţ��	���>�o� J	f�wV)�I��m��[�:i$�cEzK��~�Ѐt����C$��ku��0�r���1�2Cq(ʗ궮���}��wu��W��w�olŠ�1{�!v�0~����0,���"tk��ey�c7�DSk��U�+�>蜘M��p���8'���� ������!m�}�mƱ�|�W��Y��-,�]�b5![!p��!�]6a��X꼱���!	��~Öu�ə[��5?P�x� ��૥gc� VS|��!��B�G��i�{�,���K������]FZ�[�GGCD%��V����h��c`���;o��-aoѥ�¾�GnE��0�%,���n�?�!q�D|L�~҆� �j��CH�8�䟵��`��>�-�麥�}��K^5g��A��7��A-h�l"�Ѹ��9��LEK� ~0�o����ؿ�I����U����m(Yk,����n%Q�݆ui<,������k������C���=e�J?�z�J&q���ŒS/@��c6�=���+(� s���W����[���V탼*nt�ʪq�.�p�+���|!E'-6�f��� r9J�w��8,�z`�!֛?���*<�i�nuZ���Q��"a�aXz����ږ8j����z$9J��t��g!w���orVlbe���2�1=q���~���G�8=Kc���Q�Q�"��qp ��ԧ��h7C�5��PX+�B�A�D����M�eϢLF'�u�P��/݅���t�q�L����o�7��3�k.u�\���(�b��z��P�ؚ�,)L��3M��#�V�\b�c0����p���σ���ֈ^Z.��ުMv������A@�����wEh�3�2
+�yX�k-�`n����>8ʹ�R�� ����c��wo `E�	��knё�=�H���{7�1͈�}kU�Գ�kY݈+j�j��$T�ĳ�eN�M�E/�^�RY��CQ��$����A�W5RD>Ȟl��T��<?9:���8-4�85���Bo����WĖ��ٷ><Kaಌ�k����5hx��g"���x�X�#x�	
�����4�R�������h ,E���ӱ����f}�A�{�4����5L�D��z�7Y�郲j`�������
���b�;��س�}�����u8�H�G]BJw7�hӖ�sWs[-gb��&}�=�U�v��Y�=Wk��p:���Ĵ�"l��D�H��z�۔�3�[d�+���?�}$$�<�P��/�Ţ{�C�IB�Z��7�i��!��A�K~���1.w�2T� ��H�[{����KE��,��TIc�����j��Xȸ8-Et7�C�����L�.keV��l��%#�Eo.\�?Ir��`����V��`rr-Q\n8(�&`ǈI.��v:�?���Н�ܱ��{��961�p�y0���x"Ğ�
��Z��M�Ŝ�^�u�<�p��-`6�0����t~��z�����x�K���}MDBY4F��u"*~�|�θ���-����$ �LK&�A��;n1l�Eˋ;����o�uW��ǋ
p{Ao��G�H������z�[�286����[dKrkQ2���޸}�(�@�~���|D�y"��~Z0��'�����N8Hx���J��-��6O���b&��?TZ�5���:�h���*@8��7W��[��p�,�����?�_oB!%��#�RD%˴�^�ǜ9Pܥ4(��2�	m�s���Nވ����違'�ِ��:8����-�l[���Cź�Z�MMf}�2���r�d��K�Lp���e�F�T6��$"L"�Q�m��G�S��IݛV��)yZSG-@M񸮪��T3�f�Vo�kۂs���p�UcȀ;���R���?�ѾU<����WW��u�Q���J@���\�6��1GUNS;&����:����-^K����w�i}�N_(��Cw��@�k68�Ub��Qđeaٜ*tD�FL��#�+!���n�	�R��D70� �4��T�ի2�;"�Z?n;�0ڟ�����0w�:�	y�r-0�Fe5��B=@"La�{�����2@�M�\�q�g�6u���b'>��qq�[�7r�9ᓖ,��P猍�K��ȗf�~�~�6~�9�R��T����ޟ(��2�K�f0Dz3�V�c���ބwz�H(���-�R�����ն`X.VR��Aһ�n�=@���]Ͽ�~��D�-*G�/,��.��la�tZB�D��?u�k���;�̸8G�狙���Pq:$`������5S�f|�� X>�Va����R}5���Ej3� �'����V�s��մ�@��g7Ӆ*(B(G1�(���8"�C�yk�;�*8��a���S WT�8.$c��	��SLGu�M;�b�1�ֈ�X��H�ވ��d\vR`��"H�F��	ˣ�\�(4��X�Hi��n�ŕz�J����<W�dxW��m�ǋ�J���)jוm�e˥��o�؜1�b��t�)�����0�Q�2x,�ov��D��5Y��dpˊ	�a��^v"�N�{�WU��$�@�ʛ�R���UB��n��� ��5E7}"8��Lh3W��|>�B/���m4�Ar��#ޠ֔�����N]9Ѕ�����1"��;F�,���s���VmԒv۱N�ҵ���2�fȅH;o{�B~��W����/@`��h����݂����Xc����C�����P�`S�OF����I�$��r�EkW8L�fVgx���=2����Ё���ɸ�(�u$��~C�J�%_:�M��U ����*����*$�w��dHnk��m�Q+/b)9ֵ��q�.<��l�PI�)�%�'�P��;4�|��޾�<� X���!�L2�x�i�GA+Q!ws>t#fl��ϝ�&M7�ιY,��6XL���#��y�B-bٙo>������� [��� ���١f��
�m�+ ����nz,�G��z@���O^�/?4��V�!���.B��,��N+�8�Pn�����#��#&RB�̈́�bN�9�Nș푝�0�u��q�S=��޽|��7H<�Ʉ>6����H���@I��B[E2��X�ŵA�7(�9��~��~��~��� 9��4�m8�NL��`!�HW��0���G��^���x$)�R)ќDr�4���hU��kl�!�|Q���a�2i�U����C��v��X;����;S�v��u�TE$��������_o��t�6�������`���@�LC6������0 ���ʓf�S�pM�I�%~-q�	��J�W�Z�كS�p�F*QDDg<��.uy��Fd�T�Ar/��5|9ϭ�Ս�l����L��u9y��N13^�����*����*�1��O4Z����ԁ��n�ڈ��7^�����_���:Բc�;�a���rڄ������VTa��#=c��6��mY!���p!��4-ɝ�,�S�@�ƞ��M4'L������L��Z0�J)Q �������?��5�~���F`V~������~`;+g$�3����v^�ѕ���v;9�h��L�|S���)��;&�W�F9UU=���Lԗ��5�s����}#�X�)^d˨f���\�U����5y��e_[wc[�/٘*oJ��� �����%���f^\CU 5� �u-�9Q���U��`T���8�������VL���#<��`M�:���D$���;�s[�]b/D�o�X�z"5�PfO���a�")�Sf-��2�M�bk�`��Mx�ֲMu�f�A��C�b�����o���S��f��1OF�30B��Ep>>�Hף*����I�_|����W�hƑE����Cu�Kv�<���`�qL;��E��z�Ҍ|�{�w�o�M֤�k̗�k(\���\�C�SP�BC舑����\u�eu<y�wl0:�a��m5ot�f(LHi������{I9���.<�q3		F��{�W0��B���`QtS�?��A�����~���S�)�9��[��ʾ#m��,��-��Q������4����i����+�:�0I��HtƩ{��7�����%WЎ(��.E�Lg�PrY%X�J�� #�Ve���q"I�[��Z\��!o���b�V�=��Ο2�Y��w�9���s��Ӣ�9h=����<�h�H��a�ۊ��2�!KD=��@��v��o���G�>�g�rnN��c1Z_��m���Y-3��\o�g:0��TX�b��B�\VљO��׭)��8Z�Ѳ�FJ��84�)k�kF�K��)Rr���c�G�o�+S��Xc��Ǭ:���s�_pu�� U��
͜���d}Ǝ��a���D��z�2X�o����;P�"�[�F8a(��ذt�@r�gsk��,q甝k�5ܮ5͒���F�]���:��m(�C����*4��.��""�4�!�6}��b�o`��'n�%��_�E9�N�9�O��L���aj�ka��N�^�WV�Gr�1#��!��#^��:���(��M}n����ʉ*s��V}�aR$����z�����$!���b�A�ۀ�{x:��<X�����}���;߿�����` k{�&�W�����X#z�������9�Z�]`��5D�8�D�lAs�dKAx�,��>m�^Y� ��A�U��	��t4�Lq�Z���9��<�0.�	r�=>�8�h^���Q���8�PQ������r&����6?��,�ƫ��8ȟ���O!�S(ۼ���ϋ�����6�?�
������[����9��3�{��id�ٮ#S�o�&G���Y{����C`w� ���~�����<�\��w��j���"S���#A�B�����ӿ@��BJ'�b6��֊�&�J9;���l��?��0ɠ(yʋ�CΩ,`���k�y�s�r�BuI�b�x�&8F��B��^/2���G����[i�X)X��	^��u�xꤝt��;0��q�]>^)��b�&��z��ҠC!PL��`!H=f9��I/B�_�����[�C�A�L����f��WH�t~������.�����:������bd����>@����OF�A��-]G�!�K	Y�*���-���h�m �*��!u�X;d-�{�?����@�ѻh�zƃ�.C$�M��.���Q2
�6��h�S)P��St���G��*����3���_�2>�39��"2�("v&�K��ʸ�����w�����4����G׹�I�1��#�M��	��������L��E�����z�F�˛�%�o']&�({dP����O��,Q����� ���&�
"�}da�j��:�z��C{!��(��k�����Y����K��T� |x��i��B�����Y��*��C��~Ç :�[��D@s�_"�Η��X�3%R���TU� �3�RI5�t�拳n���]6��~]l3������b1�~u�o�r��dH�y~u��X��<���+��/W<һ�E�ٌ7��x�3��I�j��͚�s�捖Z�F:H��b��W�q��k�ENa�Q'�pn�hB�
�6�V���'�n�L�V{�N��Hڈ��wi? ��2	���� ,��ϖ�hS�v�v=-.�a*F�l�?���SX���$�Z�K������Q.��g��G�W=���A!��G���E:$J�\U�G�|~?/�y.p�����G���i�-<�R�.3�2��Z�WɅ.�ݯ�C�Y�k���ST�b_����`4-6����A���b�}���
��t���A��ف��-2�A�|�|�T��<5�'�E@������o��}M,@FHDT�|�rNAZ@O�9�U�ޣlG���U���h(P�OK��w�K{7�@t�p������_�v��{��2��ń��$�0�<���a5�:A�O�f��J�܃h8��}H� �٣�&�6#1��Z%6�&{�q��4Rv�{�g��;D�!��0:n���K6��=�<Q�ՀIR�ぱ 뫌��?��݇ ��~���)�Y����н���C�lbn�=�r�>SY��q� ��\��W0����K�4�sCBq�3s�?M�aVo�Y���c��f?��	��R�Ň_�~��� �cm+e�07�xJ���P�^�g�@	���E��L �&C�O��Ce#�*S��G���Q�Xc���^6(d䫾b�{ٚ�p[e텤 I�q�X���\zsr�o:N�8 |?�D#�|��ّ���G�A�4kA�F���x�s:���b!�hIǅ�y �2��6^���G�-���&�ռ�Y�ZI��/��U7����y;}uth`A��rq��]&Dd*�� ��Q-�%c�����=�
�D���;&�%�◌$~�$!
őK�\����PH��������\ ڪ`���5�	�}${������n�*F�"��Kƽ�]�����"0d�=y.^���I!Rdu;z�A�D�1�5�]��KJߨW̬�Ao���x���+yj�+:+d�}��mb6�Zŀ��NE`�z����tt�X�H��A�\4�s$wv�6In# j�s7�l��hL��E ��U�3�)�sˡ���x�Y�E����h��&���dv��`�<ɬ����MK�OfcER�^m�P���Qd`�.wL� ���T�v� �l�N/�[�O-۱��.��ԶҊW	��h�#���J	��;�v�3�(}Rb���{M�*����r+ނmJ���V`�gY�݇��)��6�$��L�T/ؼw	� TyI��*˕4v��9�7����s�,o�{U��X�{�9!�=�t�m}�t�+j�gQ���E?��͔��S��$��//&��cl? \*�EH�>/#���-��룱��u5�����M�医B��8O�x~�b�����{�x|dt8x��ww`������2e��?�|����R�7*�/��Cb�t��3�t1��|��`�P6��^��9��<��2y�Z �_�w0]O�|�3�K��E��W�Nu�
����U�|Y�L{M��dV���8B�ȯo���x��|�l���f�Hv���$�z�*�lmM(h���u�f)g���*�.��z��K���B�7���i��W��BH]��.{���KA�0Q8K����I�֦+S<�{�7u� �x.v��ȱ�Lle/�ӑ+J.ld#)[�	�����+*;o��%���	�@�p,2���U�f�k�u��m��RI�W�A��ey���\U�9��w�s��[�/�6�37�]a5'�m}���?%�VG��v��傋{<]l��y���#+�G�)��E������|�:��V��5f� �<��D|����)�0�	5'A;��雳�Q2ԉ݃upK����W#���Z�{ֆ�Y���|'sBbd���[�6������AI�����m"mZ@��1f2�%é�#��J�|�?�7ݒrɦ�E~�
j�,�Wc��13�R��q�h��ɚS��o��b>������P�p��!|��ۗ�Av}��U�98f���=;?H����v_N]��6�RX#�
�g�E��O�%ي,�d�A��S0�H���)S�����H���f���޾]�c���+��d��&�R����`�JJr-�E���E�=")��/n�c�*�i���g0���o�# �}B{G�Pmy�L;���N�&���`�*���ݖŒ?�K3�� ��,=2SՀZ�{��6��h�֧����E~r���Cǯ8�Txמ#�_h�Ru�I�%��q�0�I�P�r��� ��G�M"��y_J�j���Q��c��FC0rOF�e���1��ψ�����\юB7p;�CG��z���DS�� ���!�[	��;=%U9@�45je@zR�F�]�Z�b�q�M�*vQ���b�oZ�3��+��H���a>��϶�c�k��&�,�D��HD��-���-~��xX�'V�yV�|Ǽw0λW�x�$_ǝ��1qU�/�� !K��s���2�Mϊ˴U�A������b�VN������3���U�&�dK����r�����I��~O��ݸ�u0�����$;ܸ���r��Y�3?�Q�F	�!(�)8�Y�@W��I���0���W�g�k���i3�2���=@��v6v����^ϞOsh�N@��"�y4m_S��r�H��t9�2$;�}J{S�Փ�~�+���rr��I������m��B#^�gE]�q�����X�-<�J��I"�$�ۚC?�a�l�l�q�	>�R�cw�f�1i�䑿�����n�����i�n�`or��R�����p�sa7�K�6����~ݢK���iw\�s�� ]D����̱l�n�\C��Qg�H��~��rs�D0Ɯ��ƭ߻�at��Vw�����M�>tX B-�<W�d�d�CG�y��{vUA��.V{��3x�	�,�9�7$���k�0�^��Kd7�6�9q�'�xbV~$�< E[ب%j��8�����=��,��3�'qץ'l~����E�E��Hr��w9�0�u7~��f��#s���q�@ �z�RM��k�7~�l��7�z.�V{�����7QG=-Cd0�ɁR�<��H�}�f.oXu�Z��2�>7/x@|�����+%y�<FL��̘v�� yj�����`w�Q?SΨ�鼣td(��y��<F ��$A˱�(_�������#�ue�0i h���� ����ʐ� 2���CF:"(�)����ܬ'�t��Wհl�";ʒ������:�-���p���z��D����W��s�r2"UM�#�B&@^�����*���~ձ�WKF�HE��3���Q{�<8�_�EC3s�B�u���|��W �Y�{" �C�<���k4 �<��ka��9
V5PmG�E����^��_;&u��.>m�sRZx���]2p����Z�v{����o3��/	6��s�c�ʘS|��b���;,_K@ڇ�ɩ���@n�����
��`�8��u�r�ort���<f��!G-�E�N:$�j��'����yG��ȟjbAo���3�!`�K٨FooGzr�%�� zp���%\b`Ʈkm�K�WVH����.�q��p@�����jz���aAP�_���U�H9��t���~#*K{���m+���֦����HP��q?��n}����5����]um~K� H:�u�Ь�a�.���RC#��pm慯Va���;>����M�jQ⡾=��bOE�¿��V1�Gi��x�0�R>��i~O�c��������*�W�WS�.�o�k�v�&.�C]D��~��PUN��|�=0�DĞ&�7�H�o��\1-며���4�����2�}�c����0�e��Ċ@����E�%�ov=���`��̧ͻD{����-��Q��/`�lF��kyM�#���uW��� �'����A�In��m�൰�I����	�K�Z�B¦a�}]Q�.�{+��S���+������6� ��0���o|f}W_���ͦt�ߠ�čF ����!�#���`�; ���x�,E#@�ō��z�Lz������b.�=�z[����WW(M��/sl�	�P��g������y�U���J�p��S�/��V�߲�pm����ja�&��ی��r�nP�c�G��Aõp+�?���fh�$5�x_��0ۚ5�!#�Q��~ugN��~~�8g��mX�;@P/G�hG���]L�e�ī&��kw4+��€�pW_q�~�Y�٧L9����,a|/m}�ґ�p�mNV��6��@7~&�cCWE%��_M|C��p�{	[ |R�+�2(�^#�	9-'���h���hA4{��ɂ����YZq��	? �	�Z��\t�?E��![ó;F�[ܻ愀,��qT(AP�^��&S5(�ķ����W�s=��z��K�	�O:;$�sd�W5�z���t�� ���=و�'��Aʙ�sN1�Fn�Z&㶊�v��d�.��ƅ�Vc���3a��$��ťx�G<cK��}�)hA�}P�������f�����tL����-lM������F��jA5%Lj��Az��������R�����PF �٪w�X�L0���`�n��cC�����T]3?��W��o]�M�*ęi�
�$��$�����}�2����2��Lo�?9
�y�Z�5��4u������qG,����L7�"�����߮��JU�?�tޯ�m��tr�ҕW�=����V�?��͡(���Z�K0�՘]�ɩ���Q��0��w�e ����vUĤ3��0�#t4�i��W�{HA轰�\Js���c�x����cC�ʆ��b�=EAܗe�u��f(F�?��E�� �z��x6�7%V��"On����z_t-.H�|�70�g�O�́q:�O�%2��U�=�C�т~&"�^�Bo���=��1����)Cx~��n1?6�8���)+j��y�f�`G�T�-{�����=s ��ߵG��a���Q��}��F�07?�t��6$��g��Q��б��<K�Y2~u�+�^ybm��~��nq�v#��Qz�S\�m�Rr����	s�d��a50=1��n�#;	8-Q�����"�0-6`�Fv�u�!��s7c�Y���=�PO7����������9x� P&�/q�c�\圊�G��$��N^��}�t5O5!��d>��	k �O̹ j��X��c�����	�;]��r(΋$��+�#�)�*S��'چe� �����c��$:o��B^��z�a�G㽑�ع�thO�H��|�����
=�I��G��j�#qz�~J @Q�"��ݙu��M��巵R����a�����L�ze >B%8�^�W��dC���-i����Y�s�T5��zS�9j[�hr��Am�:���dP�����j��3�~��ֲ��pI���?Ƕ�t���~s!���D��n�|
�n&)��O�O����댒-�:}T�Ȇ�i��?�N��af������� ��']7|q0��釸MBܐ�A.�mTU��x��f����7�aK8ޜ���W�}��{Oi5��(�|u��²<5v#�������l��-����a5��񄛵���h$��$ Ϻ�D�~��nu�YI� ��?��c[^xz�5��SU��!J~�((y���lERYF/�}.�������;Z�X*��rb6r`�e�{�!�N�v�&�^�� �Q����_�W�V��zG���9�H6��|�f��?�W�M�ي���ym»'����q��~Nl�:�0&����Fգ�;�.:�@A�a��K�ʥ
4'Nk��LQ�Ħ=�N�Þ�J��l�I�Ɓ
�cq�����PjO�;GF�	���Qn`�Y�"R�x���F�U���~vP���/�pj�\�+�*V�	�'Ō��v�6��~9�Aq=�=�~j�O]N�B��"*F��oP8�/|���¼�*�V���Ӄ�zK�0RÊ�ġ��Č�x����>��|y6�����[�IL���4<B�K������|��-�S�����eA��0ESp�Z�dh!�`��]Ju0v�����#����}ۃ�4��_�2�VSW�XE�Yc�KA�Q��c�dA����Q�N�����!�ɸV��� �/��3U|�}ɝﬀ��d7֭-5@Sq���i"31O����� 2�1F�a��'? ux�p�:�yzk�ڢ3/$�\X�� 5/i����+�p�~��e�	!�{����%h
�}�x^�#��\/��_mҴ��[c;y&�/}��;n���	���ȝ���)f��j�M�3D�1.�Hܶ�"s�_�������!�B>���WD��CX��o��S8=��葀\^�g.2QV�i�xT'&��q]�J�8����Hd��ц��ua؜%���H�=]#��6kۂ�Dʆs9b�*�謹����_S7uQ1b���TE:�h�5�c�V2g;��i�G��#jh��K6���x����2��TA4��v\�G3F)�Vb(Re4�{bu�}�Ql���Zi$M����d���j���x�a*�M���~	@$l�&�M���;Qܔq����ks�'F�L'/��zw_�Պ��K���n{~�ے�x'�	 ��3�se*�W3��iKBD�Y�f�0j��f��Ӥ<�Ӯ�1��lE�8�\�:Qz��̺����yT,�~�ȫ�}>]�7����rb1��@��XF�z��05�GhJH�n�F���6�������X�����{��b�]�Jy/_�^n�V��hRZ��v�U�d�;�rj��Wm�n	j� 5;,L4,
�Q�
`K݇�&ń�V8�|�"�r8(A��1��:#6D0 i�Z�%��v*���PƢY��+&G6k֝��嫆��Ɨ�;���F`�-�e���c�����_��[U�Td����<#�:�G�>�.��
Y�͉Z��^d)ɭ��0U�j�`O�������Ж<~�����gKU��3���5(��果�g�,�Ɖ��J(����ϟ�X�y�u�����2�_��V�Eِ�z|���/����&�QS�a��<5L��.@�5s�����9��VZf�����rE�ǎT>c���
��U�FĦ����r������'	�:�@�hZ���6�r�a[=:���X���5!��o�'6��B��wC���߼1�2�m��y��#=>+\����U���n6�V���v�h76���	-�6
��x�Kl4}e�cj-�.p&Ň���6h���I-��/I����7�|:�Gt�-I�6 +"�}e�NG��t8�Us�/���ƨ6�����[_�[��U8�����i���}��R��7����TC�$���g�o�p2h��g�=\Y�A�x�#aݎ�� Q�T�u�	�I|[,v��]?�ÿh( �c��.� �5�3��vgd�w)EX��%=^�=��[�V��$��AX�W��C��I��k���q���w�J�8N�'����െ5�yr�G�>/�r.�ź�`��.N���H��� w���զ�N���V��������EL�gi�t�p=��&Q�'
�Y��y	"/d�Ї���Y���Z�~>��KO��_ߖ��#�.�9.��[29�8�'���g߿��v��R����p?h�tR,�NЩ������j�Ӳ��ѐ��k<֮v"�Ge�z�n������T3-:��z|Esm@*I�Iv��2)�����8���Ǹ���Ϊ��},�����cFYSO26孖������LK�� ]��1J�H	�v����
�9�Qާ����$'���m�*D99?�q�g2G��Y���p(+��C���;�+��Hc��W��@Bmurj�P��f^V�y�PY:�W~��fl�6kW���6�1v
o��(�@��4��~F��3��9�U	y�Ђ	c������%SI���5�xsX@�j��T};����F@�d''����O�&��9q3u�u]p�B���-7�GT���}A����"���2��r�i����7c��>Lm��CDe�Ĕe�3|s#�/;�y/עSQ�xT��w�>h�҉~�ku�x���e�V��]���d)�� �t�;�)��a��U;���*��=��,(xۙ��e�
�����S0��T	�}��B���3u)�f�M�(pR(���Lڜ�=]��#��њ��|�4f� \��������-!���"�"I�:�-En����H.��r�:�4?֖6�`K�u����V��_�����퐺/C��S
y��ʳ疯�>N']�����Q���R�4���˳�f�6�ӝal�����SH3R�N5�n�'��F'��n� �yy���U���V�{)^�3���|
/wK�+)ҽ�y��O�rY���r죃 ����源��5[��#ˆs��G�[	O u��&�k�Q�{�|	`�Ǭ�1�wR�{��5h�h�i��Cx�ln���n���T�3���x��F��E�},,�hdM�<<*6��L��Db���d�~�� {o��ʹow�/J�>�j��\<��O����4at�+E�1�H�p߱򿀆�q\�Q��yղ�)k��7JW��\x+��*Y
�����D�Q�j�����6p�Gh���a�1��ۈ���L��~���-^F��y����ߌl��1Lh�v	L���/�����m�C|��.�o�r�ZH��S��=�ys����=ñ"���M���=H �rF���y�Y
e��)��
)1�,7 xӒ��H�=��m���%���Iң��hO��Y�1�ϖ��D���ڗKC��Gܲĺ^"�m46�
�l��=]�Y�"�[��d2"~����3� 7/�z M��R�ƍ��fk)ZY7���3,�k�I�A��TAp@�{[pⴞPgW�sJ@�@�L�d��]#k�B�F�k��o�@Z*���Gb���^�|4�ݡ�E얹��'j<�������{]
��Ut�5�����{'}�� ���)Wyex{�&��D�3e����s�L|��< "?�X���^�(4�DR9��0p϶�I1a�Z�\q?�Lr^�&��N(�C}g��{��4�,�se�=�襮���#w��=��A4��	w�>,��Z ���%?�.�6' �E����qv�zJ."r{Z�@�q�r[��x�IEJ讌�� �2�����Ђ2\=������>��72]1�Kx��J���򧏦�n7�!;��1��� 'j�pD��3G@�c����ѥK&=Ꙕ����i�Na����&$:�9�)�9b��Q� *�ʫ�����el'lp61�����P�F�rѽ�Ӡ,8����O���{��[�P�D5u�a��c+��	^�8�ֽX�}�2	D�t�� T9|�D����U��,R�#�Ʋ�"�$�W$*��IA�`O��"��M+x-���~�֎�b�~x�����
 �|��*5W��{�mN] GFd�Q�Ӓ��
�,$|n68#8�7�F��f�;�,�Tz�E�[�sԽYf�-�&[���ê��#�����D|��=��-b�����V\�AC߲����\KW���C�m�Jc�2m�]�+�:�" 6�l	6�P�a�{�(��0�8�o=� �A˿���;����͔�·2@���&F@�Ƹ�+����(O,b:d��nC�O��f4Q�!xܥ����A?�Z���RP#�JA]f }ͬ^�����\f UQfB�(e��
BA�M�a9�Is�ԮWO�"��oGl0GFl<Ȩ'q��T�-���VX���'מz�Y,��^����J��W�~0\�:�����y}��������FT����'%@'�=��[Tz��O��w��mh�S칞���b�(�=��[�x���c+�j(~�?o�@��m�d�k�5�;�Rw$P�P%QU:��]��^A"Q�z�~LNdO��*C���C�$�d�7Jc(\?�,��FuS^�7����5MG�#9ٹy��]3�U�������B�[C�,�c� N�:"�G����K����p���p
�K{~� $��F��I5*d?	|��
�(���x�0�eqAɱ�+}P��q�<i�E-=�Eh��a}�.Am#|h*���b�fc[v:oȂ]w���m�Q
JN��]�������
�'�����h�e'�d6�X��Llqgl�Ë}�P����24���YwN���r#�a�j���IV��d�˙���x�Ÿ́��_�2�P�h�y=����d���/jn�O���$�2�vմ�x`.�л��ta1Aw���̅��S�9n�0�'�����<� g��T���h�۩�K�zDB���xSOo����{g��k��R��Ygh�_KI�:�ֶO'of�C����w9��U=�O��S'�b�HF��ѵn+�{�x��1C�[���`��
���T9�4Z#���*Җ�Z%��[�_��2+���(_�[��M�ʛ3�'��}�] �ed�,Z��S���h���H���Њd����tih�G��Ɗ��Ӹ��Syigwnf��(a�V$��#�БGn��O��G>+����]��*�� ��Y;~V�������he��e�oJ1���ǜ:h���Jo&���u)��4��\��>Ҳe�BP+�h�a>���A�P�a!;1D ï�F��Jޫü��V���h?h#�`\��7��Oy[�K�9^�PLƗ��&�+"U����s֕�����L㯪�w���Jqs��Yb�dk;�Gn�c����9�Ǿ⌏�Q���M�](�M�3/�2�f/�%8��[�͖炙��Ғk셍^l��]�z4�ܫI.����tQ5$$�p6!j�1������hN�����lc����Q�1���<(���Q��j�7��O��L�)�p��1���lR�0M�/�4/��!�An����c�E����A�G@2#��"�J��D� �R	�&�u�c���`x;�����N��C�֩v܈�ž�I�]#]�T�l���x�e���!Qo�tc�@���ć-7�&	���nTL^j6�qö��Yd� ��CBX�&�*f�����6��:FV��%�e#���+6�!6a�0rt?I�{�D�;�o`�Js(��O/�b���Y�]�3S��n�I�cO�V�MaVimY��%vψ	jV���c�#�w�X�7�9W�Vg�������fR]4Ԥ@�x��d�~kB��|Fyl�k�[D�'$��a����W@��I,<�&Ƣ��� � TT��)A;��}�`6%���#�6
�\?d ��W�����Rt�9�+v��0*��������HX�B���&��/�qw;W�b��4y'#��e��P�{ 9���XX>��<C�cP�B.xrW��Do�P�Pxƶ�������6�M�]���/Ct��旍���܁i���C�j�f\�l�}H�)�;�Lv"����$E4̐�7�Vw���Cs<���&�*�0�_	�|`Fn�;�ș�PjC�n�����5k/r��A�g�p.����v�ËV�7�o���?��j���ύ�ݷU{�ֻ��%����^s�������-������<Ӊ5%�O$�h�����FΫ1@9�'M|����|Ԋ}S>�<����@���lB��D ���l`U���|�M�ڌ�����͞>���^l`[t�D�JR�?����`{0B�y�'�u�X��B�����x�Oܤ{l!hV竔ߖ0�%����sbv��4������ؠ[%]����/�W6A�b�0!6Mn�)�t@�%�E����'�8�j��<""H�oF���!|�$5�8ʣ܋/�FD|����ty��k���$㹐(�	#�ڏ�3�'�q]�TR�Bo)'/�|O��3Lr��$�,R�=/��c��U(Q�� M�� ���U�}"e���+�u�&���)F5���cN��
c�H{��hFQl��%j/�[%=g����ؾm�	�-0��r!��\x�I�j�@���R"�����
X��S�fa�۫R'���?η�!�����f���%�&G���7�P�z<��[�RO**��D�	-/�����Ma�M��V�~��8쩕�	
����"���t���#r��2��#l<��_�
�({�ݝ%.�����f�h��\�v�si�?�7B<n�����qgg�HTmf4~U�z��:�1����\ZH|�w��d�Ǩ�oyB���sܘZ�������s�� Z�aU���Y�[jW�I�]���#��I�x�~ 9���9���=�$O!?����ɾB��(0o.��a�x�6u�f��0C:�:�L�6�P����4��f{��G��C6t?4}Q���ʘ4��p�R�|)2�}*^1�7y.-��O����)h��+1S���qw'�|`?����҂5����h��B8n0K0�v��:%�7�l���Ճp����7�^���Lv���A�_�]����=��`|�����=|�(������^S��V���hPgǱs��Ѱ"�Qzf�Ŏ��&��3�Ɲ	���Iz�+o�v���q3���D�����t҂=~��c�ї�,��C�n��E��{�;)d7�ҙ�����f�s�H�g�@�����M���=���c�JC�نp2⋐���~�2�;�GM�L�J%$<��n�4ih�n��D����~	���K�4�ݸ���T*i��b���܋k*X���F��F�b	�Z�2y%�P�&L��.�	��H�n��>��m�(���m'�����O�s�8M.�E:���-��A�h,K����o�  R5��B#��N�R����ig��p�8�����1:�� ���=���?�T��36H���^n��yQ��uu���O{���/⼎60��7J&�g�����(g%��͆R�[�0&Q�X�#�0�\���혭�g�>��+g"��/a�<N{5��f+�o�t��7��\T��G�>d[���+�\�򰑩�p��!���7c�;�4���k�A��xB�|�ͯ����(^O�^%��)gP⥹��q���<�j��6���{�����}K�Y����"+雷}ῑ�**��q�
L�����6rl[x�$<�^�I;Fb0ei�KC>���䠯`�b-��%wc��$����۟V�\ǜ�D�L6rVD��H�#��)�n����kU~|��ُZ����`6�H�u˿z�O�{�����j}�-��Mf>��?�l�}���@�`��ڤF_SC=�S�h鶘a1{V�ͯ�/� �#/�>e��]˞��b�^I�<�sv�k��$g:��R�uH�P#��k5�Cʸ��&�'�3�������L���R�EBؓ��w�p����������l�0`���m\��>�b�3��/'�e�Ա�7�tE-�(N�/j��*�ٳ�b�_n��Ĩ�R�����:�l�B�9�S`�`L�h�mw�(6�Df�Q���B���`�Zq���l��q޽+����[��9�7D�,Q�?�����\�ϾO\�UK�h�Yh�XY'6L����|��6F�:��|ⱛ�m�HJ��!�����N[^Ư/� hb�Cø��V�p� ]>+c/�[�F�����0c�d�#���B��O�l�w�ق�1��'��R�,��?^��UMr���_�R�N�J�?��a e"��� ��6����$J1�W�j,�}��4�Z!W��\qG�y#N��#0ɛ	� �j�I-F��E��J=��G�E)�U���g9�|F �����g���_���r��ɼE�
i޶v(%��7X�vuH�I��N0c9?/q�!�J:t�I�D� i��%��-�;��@`E��A��r�$-�(�2(��+��C�����Ev�YT���(G8���̒;��۬�ok1��f��v_d�8� #�?E���������n)8Z���%:��~Sp�y~�Bo�I��osH�1u�!
�<�a^u�(���k�S?��h�S�tT��N�=��ccڥ�@�gY��1���Av<�օ������Z��!;�����'�:�,B����#�(p>%����+���ѫ��!IPVo?Z��S]��|�6�2���Im�:�$�q�0[�]��h���O���<5g�7G)���9�ؠ�ͷ´m��������2������2ط|NH+�V�[��#^A�s���Ϻ�V���G�a�rK��ƥ"^	�Ŋ0��z-KX]����	�8[e��"V/R�׊����!Or�C���xp�o@�F���}����[�t���Ն��z��j�Ex]BO�h��e�0��W�c���f���%�^q���ϧ\d��@|4ht�`cT��U),}pQ-&L=�8��Q�h��<<��ִ�7���%coXz�}����`'pH�ȋS5�f-����`R���Խ�g�H}l����^���K�a%�~��߸%��L��iKج�	�Bҋ`:�-�����؋�~ϚuB^Z0�δ�ES�����z�5�r���
��|jz׿��']f>� ߄�s�WF�1ST]v	a[RI`aY���-�|]Kl��{0Ht|�)l�ؕh���y�
ς��8��:�
PrkpbQ"G���&\�δ{9���a��[�f`�H`;wJǯ����=�0V���u��M�MY�.��Ŝp�*��gS���g3XofϘ�(�I��'���y@��~�IK�m7�-��x��:ŭ��:�ʹ�x�Z6�kI���[�7�r��V�,sM(�߀[vQ�����vyb[���@�\t^]�-�� �w�c���[���9�8�oR�.�X����:�[��<2n�����=����Z0���|&�n/����M�8�W�$B���Ab�v����|�"[N@�x%����m�,�h���oTLz���Җ�KCPc%zwΆӒ�oZ6�~'�".R ���1sW��kxC.vί��Ǥ��v��ƹ�t�p����
��ݕE9���>�z�!�22)AUP_���\��R��^ۘX��]p����O@�L2����f�JF���{�s2D�U�E:�+#)ml��&x2=�ՍSM3�q���}��-�������З�(�*_]�1�Zpu��G���;���כ���2��O!:Zdɀ=��ù�*�*'�;�<�[�$���~v����Dr,ƫ�K�vx2�#�Nuo�}�~=��{�^��c#%W"��L�E���,���	a	��O�+�-�)�pC���-wb�+��8��:D�'N�\@�������
?١��^�����E �,��]�eG�=k.���	f�����h7
���`S��K*����P^$�)�W:����`P��՚V�e��$0_�b~
G�{��u-�F�;݉� �{th�x2��l���}�~[�3y��~˹OI��~��D��P��aTI�y�K/eS��@PU�?�� Sq
y�f�{QFF�C4Z~v��0�E�<�C����噄[��m�MO���t�Zޮ�FZ^��Rx'V-�*�ףz�����/�H�I�uql���a.�a-���7ص�d5���QǕZ��o�4ndU��P�ޙ�K�
15E�tꃻ�8��-:��	�D��y<k����)�_������Y���;]��J6���w���=�����kI{rǆ�}+��3S5�K�3n�:r�	�{�����A���f��_���\����{)J�Χx?�����X�D�%�k�>Ȅ��	�����kRx�3�@�	��ȺN��
����<��|��&�0x�.3,��B��xe(C�Ro
a :b��,��]�6�i]�颶�~|a{W�?Њ�ɾ=�f�?�^�\u��<����z�\�A��綐A����v��0�x�UȩсP�B�C�bR�p�����%��~��v��3�a���l\JY�i�>N |�S��gjP�\��4$8@�;B����'}R�U�+\#�Nsis�Y"���X���FDY�w,�Pll�0��p�u�d�?��u`�S�oq �S[�,�8;�4GR@$t����wӔ�ʻ�x��G�;m��޽w=y}'�C+�L%vu��CU��j^�o�Epar��b��ɦ��n��b� /�������X�Br�T� uw�Zhy�PO}��������A	����IW�ە�ߴ�|�#w�Z�3��V'3��C%�]��!�?!(�d�����E�YY ���]O$���v���.b��������3����!!�JR��3s>���5�ℵ���$���ۇ�oljnw�8PL�QǷ���};�YE��h�ՑX;�Tn��3��f�=�a�d5m0a���Fo��>��)�� �EF�\��x
�.��y�_W	��ђi�*Dȅjq��h3l<R9m<�J���p��Q����P��2�T6_���ko�9���[A��N�O�F�2X�k ,���41��+�	�zmͲy�
��4��1������f�2��d����-���|l����߱�����"AX%���w1wڲľz�+��6��4bv4����E�")�zs�Uc�z�Of��������d���$����	��נ�#B	f��r��ߠ��n�@o����Ly�(�%�oVWޫ9�d���Mh�Phd<��q��kH��5R�����M��Yy���D��{�|�t��:�MZ�����Z���{zHS�UE�\Y�������7��cg��;�8�I��	�(}G�Gb��ӑ�fo,����Aɀ�f���&�:2�m=(Z ���r���@�L/����2��&�ijE#�Ѿ��z�v�c�u�M�*g׺��:;���I&_҅"�'�!�;/���
^�=%�EbI��]O�+�p�>�,J`�����,c�#� G0��̫�ڷ�C}�B@�(�4ׄE�E�C�bN�Ϧ��l���ϯ�9ϫ�{�	��$K��5��E��h�ƫ&$xU8�+��ekJ�(��\J���_�1Dvي��� ~_b��p`���G\<�a�_M0��ו��w�C�����9��a���*|J�+^�	��*?C��gO�B���_�����-M�v�����@M��[a���R�g�u�gm�Ơ�2�ţ&�G�6��{i3�$e��I�o(	~����x`U���s�:���u�a��XKBI�FI�+?�Y�bF(�>��-�KAP*����z��F��g)�W1 �x�/�1��D� +�%.�a��D�������25O����0s$1\A@?l��mp��}c�t(�����TԜ�_��ϕ��>�:����<�=�2t�B�.3/' q�k ��1�й-H��8���Q��݌j�h��R|�d�VngWű� ��f�-׉sFD$&��_��o����~9��Q"�V��8P��9�ɯ@Ԥ��W�>H4
��k}6<?�X��,��%*|[<�s� �m+�6r]�Z=�����᜶�Y�c1�+��dv��y��ZY��r7�su�V�,�X�iV��V0���}z^j�`���cO�0���x�1�v��i������+�������z�?��/؋�KT���l��$���|ɖ��:a�?ե�䛧ȳ�@�J6 �����`�b�6�A}�p�4��+��)<�G��F�@7+eυ����G^����"N��H�p���L߻\���x	��!���^��]���؛=�&`5�Y�a��g`!�_�?&Zc1��^͛��ڟ�،����/jdA��5L^�R���]���o��E��j�Oi���������]��A�k��=����7���+�ly�����O�|X�˚���e{&�i~`X�G��91������J�v��n>\��T��Sw���#�.y:�C�2~�������Hd�e�aE6���K�?�8�x�g��~I��{7��r�8J����Ux���|>�IM�ꉉ_���2+l֨m�,m�A�欁��~�/?�W>%c}��+�Z2�������#����D�W�4RoK;��u�����zf
qZ 'Q�% ���\�s��� k��[�v`I�&�t@.��)�cWy`
B6G�y�a�?ufSnğa6�8��cT|27ԍ�\x�`���,���6��K���=Okŷ�����m���j��� ���i�"��%7��T<O�i!�������CW��Ne�&� N��� �ә��dgࡹ��.�WXc�Wl������e#�N"B���\��t���ߢ��� ��BO�)C������n��|����G*��0f) b`��顔�I�H��^���B-�X���{O@�bI��mp��R됈���y��D�`�HS%���(o���}��+��%�E5��������w��jwn�ViIq���g���K*:hq1��n������!krg���^��̛8�q>�{�y���Ґ�;�@�W�)/*�7d�vCliw���Δ*K�;���a��������Cb���F��`ӕ�;ث����K�P�q�ޜu��I��m(-�گV��XE��j��&��)������@�(��i��� s�7�yjk��BF�ڛ
�9�?��d��;d)ɪicPc��������:�l��t	n<��b�脝�:�T�1K5v˗V*ʛ���EOXӦ�YԀ ��Qq�uK̸m�RN��
����=A[�t�딸�i�u�D|�0�"L����$IS��\V&�*���[mࣔ[�W
Y�R؄��S]�1��>�6�zJ\�����(��F��U�c�_y�q��,b/���s�L��GOw�޹䲨����.��1����� a�ۑ�~�#�������A5��N�J����J�K]��B�:�t��7PT���G�V㯠3m���e@�>ɰ0Um~�j�����?V�7�]�:���bե���F�ǐ#١��˴^�g��N.?̯����vJ$����K�;s�N#м9
M��;��	���L�g���8�"��Mds�	�����2���n��[8cdAm�Sjy�Ò�~�l����lnE�e��k��s���&D�Ҩw�Jk+��a���r[�IЀ+@��T)lq��<.�e�)1�,��!/��WJB'�N� �
f�n�1�k����sw�1a��kA���#^�L��!��X��y	h�[/��E�ni������,���w	��G���_C�X�+�	Q}#`�Oe��e\�{XXqՠ?�ٍ)����$�v鰺q�1QFK��^���?�c�RE�V�=��D
/�n�ع僓��A�b��_q[�`ˇ���6����d�	'�M���nc��+��d`�V)����'�ϜW+�6|E4�����b��1����vN�;T��~�e�9H��Yɸ�+���毑���O=A�)=�H����MHnĈ�+QB_��Tp�f�^�4�9�����s�w� Ƌ�㗈������ H�E2m�_&+Z�쓕�+��������,����Hk��!��p4J[��X}+^q��3͐k=( �2D��
��� �2��?���؇Y��jr��|[1P����x�c5�S�Z�
k�}ecC0�����x�2߲�^2��ex�z�}���u0wf�כ}T���B�>1�qE}���e�L�g���W9�>��k-"����a-l��FG�<�F��gZSbE*�_*V��a���n�O�0#�)p(�f��=��DH�#sF��L��[��=���(�;G����yb��sڼw�n��U}i٩��3��Ӥa�-'�R����k}��Lp�-��t�CM�w&������G����hs�g�߻�+j1���
\����:f��.�)<�!Ҽ'p:MS	��j�mB��#`��y��d��B�%��ܛ�r���3���w�e�Tةxp!�<��[u(`�ϙ�6��Ő�֎"A��P�l���V��L.�<5�j�j���W�=�3�.�uZ�.5�jk���?@ǖ2�Ȕ��8��x$�<r�P��Z���p���Lj�	cE���b��:dݙ�EM�e.k[#^��hz�s�+i�-<��ʰ#�ȋbǈ/��[l�U�Q�Bf�H��S\���UV��~��.����y�b���*w������Չ�X�m�g�j6�]�m�۽,JG��Zϥr�����T�˵��:�`��=�wʟ�kt�a68�e�Gp�+4��kz�B�؞��0�jx�ja��ܾ�_��'b��:'�Mm�s=m%є8�=M��G�Y7Aa�{�~(������ ���I�q�auSq��߄I0�@�˼����З����B��W~�rn;�]�\��^�c��J���2��h�:���#D��AW���m:m\�#��6�uc�"�P��N-6�#t)-�J��<)��zj��b��j}�e~w��\[��0q�/�����Kh%X]_r~(�5Tq�i�!�^�����WA|`��߂l����������@?e����1Q�}E�3�סF�uC^�O�G����~p�A����
<����;D�lM��a�^��)�~�+n��=hrz�EIe�'�P S�`K�drl��w��6H3��	�"韏[����6Y����6�lFkb�W��x�� +��-� �i~I�o¾@��&�RY�]P�E�b&L"���IpPm�ߪ�5�z����6v=V�#�?�������:��
j]0;�L��]3-i�o���cqk7��JN�����,�����vu�KO;������(t�5���+B`zTٌMr��ڂ3�ST��J8�˦�C4��Z�k�P*h�ݜ�6+����B�Z����[co(!4�`\�t�q
��.�"�plO�q�\0�-��2[ �=�`�Ϳ�o.ʎ���?�\$~�13Cj�0iU��؁)*�G=a�REc?�c�n(�U}Q��5Ë�w��p�i\���'~[�3B���L:�3��W��]0��Ì�i�-�����Z�]��Jf�J��/�36R���+g�/~�Z��� ���v�����zf��1C34���gus�f-�ZZ�zxٔ w��k�j�F�u.��
8u��z>$�.L����4�5�>�Ǐ,�B�c4��#�h��H^h��zAKq]/+�t_��֖���:�L�m�^�1���d�.Y"��������#�%��|ӿ�p��9���������A�~�F�D��uG�Y1�Vi��"�;�����k�vȒ�n��I#7��~cD܃�f5ڞk�>�\'��yB	oZJj�(��O�m��|�rK�Nw���i!㚿r�H��*i��"a4�����c��d�"�{�6v\\�6�6-�P�z��$�R��f���Ee	��`b�u����y�:��޳\�(X�L5>��J�CFh����֥"���Q�n���P�AB�1�����BĤI�Q�-�q��AI�d�ys]��1��(C�m��%�b��|Y���k����2����R���W>�gn*)�isY�6%;�^��6a2�OT�"�tbeȗ�&Z�J���+u�D��Ĉ�� ��d�z��N��A}uR!�N�Rb�6(��o^��3����)�B�[�y�7��� RXv��b�U��H7C�CB�{n�d�v��}����5���t_�fgu˪�"�A'�Z��/���,�mʒ�������vs)S�@�
R��C^��<D��`���;��d�4TV��k��,��������j��g��+�f-��&Q@9�6�H5]�|��r3����U�\#Y�¢a�B�l���BxХ,�qtb�%ӺR
B3,M����n!�4h>�j��!����
H�k�!�(d�K��"\^�{{�\��10re����E&!I�۞��䟲� ���;hm$���c�A'�ŐZ�c.&Ň^�~���[�[2�5��Ȋ���	�����pgsB��M�%A8��SU d�.��^:{��8t0�֐��)��Lq��;8J���}�Ǔ$*w��'e���
�>�d�<�d���YJHG���{�+������A�E��]~r6>ӆS����0��b7��d�ĪF!,��/4i��q?�X��˯���[�N��/��4�����눘ĄRF|�(8dlG__����ѵw�<:��nO��
�%i�$����vaT��d�lb����W��_���o6'��hM#��TM;�%`H�B)5����xP>��m>�l�o�&��"~�՗E;����ӄB��]�waP9�,��ɱB�W#F���Gs��)G������;v�oN�'������j`#m��Q����@OLa�^��ԥ
��Ќ{�@A�D�H�\K���>�N�r'rI��i�[�Ln�J�e�؊VM��������$7��رz̿+�E��[�웖4ƒ�y<�dGaa<����;�v�G��ԭfn^��2�GD;1藣�D%$°�O���Ϊ=9���vU�wqRl�8�S?�#T�n��2�oD��h�z��w^��v�2d�F;@Q�0��j��I�u|����>�Oo�r�O�8��9�lZ #���8�8o_9�!Ҁ��/6#��>��Y�@�Fv���x�+D,�����vK�R��g��K�lz�`�l⠚���?AH�(�����K���l���l�D���P���P�Q
)�+�aE;"��q��y?�q"1	t�0\?�vL M���zb�R��Ûǧn�YٓKZ��\�_@,M߈>��s��2P��Ñ���ǃE䕩���[�c�8Y�������~�C��/o$F�@��^O�yM�8�kP��qZ�/G�=��)�B��)��oۦH���R�> nF�K������8�IO��E5�-�E�`�*[IPY�*�iE��3���Hw_�V{I�ч!�g=Դ�����gS	Z����V�8���9���n�����{�]c�����b�%]86z��*_���;��p��C�W��>'�'���цZը��H�Zr�ε;.f����\���Y���!�p=i��N��l�M�pQ�DfqÀI7Q��^���s%Ϋ�����EB�kİ�C�<Dt�|uv����J�R9�9J�6�s]�էbmrC��t��ӣBL��K#=�HAw��@��#�V/����N���j .�/7�p��.����ǈ!U��Tp�E$����	'L4����k}�(]K^b������ʼ���AJ���9��6BJI�����2"::('�f�J�Pa�\�ge�<tw���!�C����0Rb�Q�ʈ��
����[�.K�ѻ�^�+8wl��.��8����"����jb�[�F�Q}�;�h���(��3&-P����
������q��:�袉h����� �x/,��u�#6'�[�(����ur�]{�����~#@�P��?8�оZh��[X��ŧl��D{g.^��+J\�7�y�8�����%���3�w�����9�Xts�1�O���pڈ�Zz�!<"4��~igf؏�wWn�[�� 8Sة�K~�w���'�/B 
�����}#�$CB K�邊�EY��*S�����Z�<���#L��`�n(�j��9�:�?��(t�I+���C�1��'�K�J<N`H��2��њf����<�m������+<����?��������v�˷���\l��7R
��:� g�|���P˯���7� ��*��@������\۵��&��R���oM��lѽ�/1��;2=g�#�KU䠲�ֲ�<����Nb�m�N��o3{����y[�����xq%�ϐK���>O|���a��h(Ӆoޘ�)-���0��o��-���'��6����np�F��������Qib��NKJ�~�&�X�#(p;_[����\52��*��g��&���ߴ{��2a0���Q Ys]퀭��:��n�\�eG��9�%r���/�6؞>�"Mo���� ��}��V<��}��H�m4��.jlÀy�x�,�x��2 �����8���O`M���M�~�S�M��<�H��v�Pn�R�$�+j���X �s9�Nu�ϩ�x���f����������6$\v�V�_��mQ|�gċ��
S����I����2�����W�}[�c�E�`T���[�f��+P����<0�Q9�kI�S}C>ߪt��Id�rzI���xUAk�}B����XS;y����xD�&G3��g��U�^O#�~~h��H+ ԯ?@����'�ܥ��+4َ�C;|�h[���(b��Ab�b�C���䨐o�����aH���f�*g"�qǐ�z�������$l���6�g�Q�w򅔓�M���i&�^\5[}��R��A$��o@?{��f�� ��&��T �>B�\�e�R���h �f���`�c1��I�3`�eл�f�Ȉ�m��������6F�����n���0���oJ"c�MP�F�#����L%�S�kG0/������blKK�޴\AiP)�Я��!1��l	�3/v]�YQ���d9�R7Ĉ��" �����z@����.�h\w_�7a���ȝ�"�\wlUg�����Y#�3��Ю��ڧ�T������0C93���.��iZC��ޘeV/���V�펓�N�N������}��]��f*)���8MN�4�j��8Um� �	M��ATiZ�:��a�jςSA�N�b�I���j��cw���(�C0 ����/�e��\��Y��3:���'��\lN�P,�ɳ�~�Q|���I�T���,�v�;@�4P�r�MD[ґ��M�1�t�K�B2.8`?ԁ���!�kB僌1ݠ��2��q�����djz�"fX+AY�r`�<��K�;%#>2م�Y�r;�ON$�uO�:E�=�^Eb�bj����k�M�`�Wz/o�L�9�mB�& �e3��#$��sN��n��|S|Ur����F��� Y���N���Pu}�H7)[ϔF�9W�Ő]�2�]��6-�}��q����)�`u� �����s"�INX���d�`_�:��rWL��,T�֙�uwac������a�b�Lh^ܽpJY��ySx��Rjp$&���-C����m)D�@"�A���Ce��['I���ȃÓ���+�Q��@n��ר@�<�ۣ�O�=��W��R;	�(��A�~1ݕ�7*u�L��ʩ8�#X�]�5�Ă��_-F��Ӭ�@���tV�b\�`~��DO|����l[3k�d/���#�M�U0W.��p�ܯ�j�k#�,� ��c�(���%<A�u���ʚ�#��Ǚ6��6t>I��y����/4�q�d�$��2�,�����Xd���Q7�ݏ��ਃdE���X�M�5�A�f�*W���v��!�n/Hy�R�R |��7
E�eV�rD��h�Jf�=�H6vX���ў��!�2���گ>�u�u@�g�;qӔ<б{��71����MBV����Tf��<!|����Q� � �H��ᡅ}��G;�SVf��S��M�B(`-��4H�%@v�9u@U����)�tJ�Ȉ;x&O��ɾx��bK�v�?nF^�C�s�	2S󐵖+�Ep�J �H,�X�OJǳ��w]^��{�f���v��y�؇����m�=�nnf���_~���\)I܋5��	�ǗG����?c9�b�vjV.�F��0�UC�7H_������4]̲����\ڝ���u��07����^���?�b�]��� ���ݒ��@�U�Z�[��afx7��� T�=zے{�i	�����k�%��@�z�Я���\�/�m��k!���A*)�HM�A�fMY_x���s;ҭ��7O�aA�G��+[G�B����|汥Jp.�l��`����G��5Nܝ�"�K������:[+�{pw�U�M+hKP�۶qP��)�chG.!���U���
��n�ả����~oQX!J˼�R�~�b�E?-&����ޫ�S����E޸'
�a�Y5����o{a��r�H۸�.8��$V�_D�Z�1�7;����؆�Ok�3j�@�Y�:~Sd�"-��GY�a�0�&Q�6��C���xxD��SLΗ����]k�&���Q7�ΞV�i3��g�C���g����|���pf��K��x�z�'��Λ.H�*2^nx��Plg�w���,c� �Yp&�k>�%��|.�'��~N=b�Z�ـ:hs�0������{�pT�_Xn�6L�#z{�T$$�bJ��{u�-+9ē�x�`�b�X�<���+�u�+S�ٶ�4���N����iϙ���i���h�It���^Ĕؖ�":�wq�K/k�+�d'�#f:6L]}~�:��#���ΓbNǎ
���F��;8��G_ "�������Cq��������eh�,ѥ����G�	2=^����%q �W�{��[ƀyX���H���;&Z�@�\o뚴���U��N�5�OX� �̰M3�U���I�3�]!�i��.K���53�v�v��d�3����Q�G\;K�������@�`/{o�,P<���}���+{mn՘�{����+Z�+���B(x�О���i^���wWr`��٫%����\�Ļ��8�6�.:�������6��=9�"D ه}�ӱ���ߗݑu~�%z�;��B�1e"1qh'(!ιy���縤�v�I��!C����p��s�Z)��S���ZPj��&2"���������+�ḃ��wֈ����9��%�h`���gT��7��C�� ��;�-���^R�t�2�!��0 #^�7V"�Ь���qn��s�ؖ���u�,�����c�o,�)��E�u�)5�v�D؏uΓ�8�����(���{)n�n�g|S��K�؁E�����Q�V�ߔS	���~0܆7�0w���-FX'��q��@X�:Ij6<��\JB�w��x�m��bo��Ǎ3Ssd�6U�9KnŹC(΀�˕c>_�b���-��䳋��-��O?C ��Ⲉd}^*3|��NU������F�<�`/)'�*�`$�=X��ܿ3���߯�?�Ʌ6�����DU+4��z���;��wBev<�O�S�g�i|��X=eH�"O��7��4��;��u��Gy'�'N,/8$���(�*��3���4q�ntO]���f�����������v%Z\j̜~&�׋�� ��%�0"ա{J$4�ź� ���1S�褗��>�!�ʫ��Y
e-]�9GZ�2��F뻣�E��ff�
j����)��^�#�|�}#� �˙f6)'˓R�J��T�x�������;U\/F<i��j�̄h ��q��Yb/�}ǎ'���1A�=������<�L�e\LXC^�
+?�_��!�Hi��3��A��I���JD��f]��2���1��oѿe�]p�\�@����{��JJ=Z���,s��0��р�.g:�u�@ax��Nfڼ)�(��_z����@����z<.�Ҙ�j����,a��b%8�'��X�Ć��!� X�JE�J�屺�$�?5����#_�'ڪEL)�;����<�.�x��xE��RK�p��7Y
��k'F�]���t|�t��dI��#�����D
���a��yi��a���-!�Pל�eQ'���U�6�'h+3;sCˬN�W�@�-<��8I���
�_W�a�����ï\��#�J��wEI*Г���j�6ʘv���'�fw�.�t4۴P}mR�d��N�h�Y
�1����C�Me�D���fq�Zǌ��+�*�o�E8s�9�n��h��D;1+�w��s�w��B������>;�4OO
ʎ�W���Ku�wC�:0{Xj���/�.5EV��}�jp�jN.��q���o�|d
Mԉ��n�=XE����.�>��`%�e:�>Y�� XB�BVb�g˂��G�)K50��+���A��u5�e�#�"�b����_�� $�����Yy�O��N���4����nu����Y!�g��1��޼0�-jKV �J����z/���m�	-���5�f�뱀B��=���\Bi���-�d���Ttwz�;Hj�Sߌ�i����<ߖ���)�}DσmDA'������N=HI���(�����:����R�'kp�ï����������\S�SW�Ǆ� ���Jk��n�DD�{*�=Y����Lˮ�-`�ʒa�o�d��{ua^��M�Pn������S���B�CX�y�=&i(�Rq�OAI@��h���H���5\�FP���h��h�U��\*8�L<[��uS��=��wf�wv���N�����o�@P �u�ǀ�vb J����S�mC���#�}}!m�^X� ؜U�ٮr�<���</����=�8���w2���ɀZ��$*�EXM�X��/�9Ǘ�cgSzXܲqʠ��|89%\��L� �oe4ϸ�*Y�DC�5����k�u �&�_���2�,��8���a;� �w���@h"'our�RB���'$DӸ��此�Jo��,��}v=�'
!��vB��3�B��ǁ��%��+!\r���K�NR�(���y�@�"�;��̐�~��%�q�ا�M*2���ߏ��񫷾���w���/��&�T�K��"�t%��a�V"��E��bp;.�4�f��/��s�N�k�gα��>�j���!�R������[]ev�W'j���(�x�	KP�h����h=��"��
�)��H��,]z畍p[E��!i׷
�
sE� k�f���z��z�7���@}mPm0�`@Z��Fl?�{�=��݀zK�q����¾F��ר����Ŋ�3���J�:��,����c��Bs��ԵG����P!ۯ��+
��f�����9X��A	��aZ������|���o�1��%�hP�C�e���D���[Lݰ\�J�b��"���/��;�����r�bl����Y����ѹ�CD[�@\{�fI��'O#�ö�OE�x�,��<h7��9Vt�}��U��5����<�k�d�6�H�Gƻ�\��WJ��0��LDw��M�^X��Cỹ���@��>��!��Z�?��S QK���Zn��b������5&=�~9�X�`�m0�G����s!���ߞ���~���3���W�Ax��y�2F��I)oF�f/T5�́VE���^Ҏ�9�d3~˜_�o=�=�2�3;�}Y�UY�����NF>[���kUZ�E�q��Y���ݴ���t�������M���,�7;f�Q��(���߅�gA3ٗa�I��M@r&_�/���7��IQ����� �j_0�9}���^a�H�%�H��	V�3������x�H������	��t�_��=j~�m%~"(��@3�Lw�����\����Ǳg�!��,c�
���S|t(Q�uP3Wyȣ[_ru�Z9p#s���B9�{ÛAJ�i;�J_����|��Wݕ+���X"]J����LB�B|��i���'i���_�/2� K��0���>��p-��E�(z�Y�僱J�Rs�#�C�f_��lQ	�j��� x�k,u}\�wd6���
˲���TQ։�6��tAh5v&4?�	F|�V�H�<G�O}M�E��dͅV$����H��ڣ?Ϡ�pE��&��]r�>LB�𘠽əyu:Scl���Ll��ꐰ�{�HCu��ޒꍏ�k_����	ȗ�K�#E��t{M:�B�".t���: �Fo��?Lz��~���ͤ=��ҹ4��>�1=1!{���9�|`a�ʆ�t��
��a��S�v����$]}[H�����{n���-|�"6`� �\���VܧG�$�O"�)3�[���.��̢�#���v�6�mU��I�)�ƖjD�DD"�{t�F<B *�Q�)>T)�m��/7����=+�����qQ|q!�ע�EGg$߰A��l�m3��L�A�8)]!���DS�1�0 �
��
�.Y�r �R��V��"�����8���)��q���=�J�j�����-���I��M���IuK��V��ПV�.zlf�^?s��4n7���ry{?�ʆ!�X|���0X�$���X�:O�Ⱦ��tN΢1`��V�]���}��nu�[&G	��홮��k,�:fr&��\�� 3�K�� 	�?=JD!�R�H�>:Ggdg4Smi�[���A�(���Qq:�����-����9����2L��.���E�'����O%e��� �Eل'�FW;,������vq|���&�9�I�l�s��>�1{�E"��$����5]�g�D���O\Z�v��	�6J��mC���ѻ��{ɨ�o}O��3a�p��(�i�g�L����w��@�G�[�F���c��|6�<���V6�#(����M5�`�9�I���CeG�4/dg�\�ϕ�T�ث��*1Q�zb�,t�MK�T�e��}/���s�ʧ�����[����VI�����!�F�^�I���z� Ү�y�6��F��Q;��[�mԛ�	ڽ�H�d�k�Z���]������{
3�����:����{�0h������(n5$��l.�ǘ���Uʌ�����2(%6�cr���wٟZlq����-�1v�=,4#���*�~\o:��Z��$�he+�8�C�/]a8,���k�����d��z���h�X�b-�=������%��Pv/��wʾ��&N'Ž?Qm�4f�4@K8*��yOQ�o1b�J`�\`����ɤ��.-B�;�����J\�#��jH���������XD����,얅k"�&d�[��=V�R�?f0�?�ԘNE��l�qfh�|.�壘c2���8ߵAW��Mg���J'����Fd������� �uV�;�g�H_GX�m��cM��iYm!f���gL��."O,ߩ�S ȥ�_���G����-"��g�U��.��Ə���#o2G�}m�~�Z�+O%<�C�J#k{������^0]�OJ��1�k�SS���m�A@�����/.�V��%�`��~�II�<!�^�jp��OL�s��|�+H��mk��3M���r��Ҽ�\PIyuT�͝��U����eģ�e�wR��2�
�\N��j��%���l� (�Ӄ|�Wkh��;�Q��`9�Lb��3j�s"�an��V����[��;YZ��(�hN���QOyvO{X3��mdw����8�*� �TS�����Uk`9���,򍛐p�c�@����7Jsp�
Q�4���=*����!�~���1{���[V���V�2Ν��2wj҄h�z+#Α([Q��kGy4[�8�{r����CWI�I���V���d�u�UՎ�Ѽ�iU}`<���V.���V�=�����*=?N(:��/���U��V��{2���y�ɝU��ﷀ��i���EɄV��a.�������n��d6e4(�XbC�O��c/�*H^�ҝ����gP�*�=�6E�ubSO'�N�.-vm�ki��!2�x�ō���6��+؍N��N�����$h��NZ�u�pX���M^�`<	@��� hj	���lb�� ��s(]����F�f?G�)Nm��_+���d�4�
���b��Y�hi緕���t�)5�%8���ҷ0Տ��.mY�����XβT.Pͻ���?G�j���G"c�Ui����
)��n@�]���Ë4,-sx��9�ǖ�"���6t����-�=�Q[x����C��6_�j�H��NE0`�&�4��N&�X� ~�a��Jh�� ��~����kż�ZY��ji�!�9��/� 66��A_�%�+Ĕx?�b
?�����´vF��\{�J��L��^w��VI�ef��~�E�~Q����`�*ɏ=0	�<��gu�8�3���#_X=.��*�[��!�iƶk���2��[��7{>� NjUrI��,Z!�|Y%]�I�]��Fɿ�c_��YB�
�c��kDlb툅�� >zL4�k�"T��~hs_1?�� w����)�6��h�һߘE��D��O5�5-��PC���r�vʁbl�[њ��,Xu���
V8d%A���X��~G!�4PN4~��DBI�zN�PB}���g^�q����l8ä!�>*Ue'A}���^���j�M@km����ET�����R���|�)���?�-3�-��@�!�bT�!>	��gF4� �EK�iY*l��A�lZ68����*��\���%�S�>�'�g�&�>�*�S�y ���bU���UE�]�":p���	�T�2���u9�+ ]BﾞJ�0%�����
��GoU����!�+cz���:�]�E R��8.�b�*v�|>u&e�7.��wL���>\���M6��L_緰T�4uQ�c�3k;��vap���a�=�BNP�p�,��)Ūn=$�H9���T��d��0ˬ���<�a ��l��ܯH3r�D9��ƨ��L>����Y���WՒnp����C��}M�&�,��,9Q[�5����"�ۏ���C��(:����B>Ȳ���~�>i����|��4�3V�
[+:�5̿�O��2����w2{H��=�fW@��9ʲ4ˎ)$5E��5%�:b���@6����mr�I���P�sv�S;���%R�'X;y� >��;��X�kQvx=3K`Wi)=`�n�]1�tB������n��"%�J��,5�rtҏc�H�:���'`�2���`��w�9��iƣ��@�.�spl��S85q7x2^��������p����,�
rQ���Y�l{ՍsY�Tg���߇��^1�s�ǔ�>�����CNVC��èA�����\�L��@��Т~��0yBxv��������vע�f[��ey�F;�d��B<HA���(�����a����;;d�r�1v$�'����ׅ�Q��;� ��DY@~x�hC<*���,(��Τ��#�;}Û$ƾ��j{����
�.ءs��p�;t�)j������v$��epz��.zv�����+�$呒u�{��Z�"�� PM��i^%���A��<�Ѕ_ɰKer8�Lx�3Z�
ah�1����&�K��C����6��0�E����ʝ�ٲ3C��B�V~��Js~��#b��=��s�ֽ���xc��ω׵��]�H2��տi��ds��qO�|�X�u��9�4S����%��PM�2�K�њDl��T>�	�0���q�L�,�޹#W�=���[U��٢�Yl Cu�X
icJxR-3����.U97���F�v�g;��[x%��:!�X�"�z����I.:c�/�^i���;B������ji�E���@�#�ՉӛW���Y�����z��hԑ\ 0�W����VnR8�NT�0�Nl$"���������GdR�G߽�X��T>�M����_Y�P�b��=����:گ�:J�����x�#���4�>��s$�"�\
"X\������9���+�hpg�:f��ۚ[ǟ�����%�c{�t�C2-N� N��Ѵ�M��z�4�����Z&+���4ܮ^rȈw	~n ��)ȁa�mC�@�:Kf7G�Q�����QCqE �7p����x��#������j�MC���a�8�Qp��.$/u8XX�9'�Y���B�����&�)��#����p������,�G_��s &�;;�T�5g땖V�*��C����h<5M�~6��&��&R���u�p��v���(�\q��'ώ�;�dz5��_�y�]�V\>��=JV�J-VaG�G+(�v��9N�r�"'?O�]� L�Px���.p"���4΃��t$��F�l�_\��������ŨYytF+�����M�H@Ue��̱eY�Y��%���`��9v�����ҟ絧��x?D8I�{%� �+ΌR4A���S������c��Rw!I31�G��$�&z�x�]�^ᑃ�N��vi�k�#_�&�������11����^�G\��w�����4��0�N��a��"�4��R��B`%'s`u�n�	j�kW�(������aF���6OYX�Z�(�炶�>A�Wp�H�ˣ�����Y�?�6gZ�O��]z=�f��%�"E-'�u&ql�Γg]����ȸ�g����Y4̻[��t?�cb��a��be�68��|
}���}n�h�ġ����hЧE�-���a!��~6��� W&�e���q5�zA�_�؇���SV�!]��E��|JGl�4��ѧ�^p�'h��m�fǗڌ%��Z������@����2�r ��;l$���j�v��D���jvx[Q韹Xj!"�}��Mp��aRDޝ�yo�i%
���>[�)G8ؽ��T���2V���2t��X���.��%鉩��:6bf��/L�1��0���}?sc��S��ݤZb���j+4j�Uʃq��B��e܍�>Ō3�~_�L�vߕ�'�_�����|��zq�1��fGߘ)D�}��ڧ�J�=���˵ܼ���p)yt��s�"��g�N/-�Y�,�-IzK�m:40l7���ݦ_�J��I��7�/A�(	^�-/���,t����RW˸�0lU��˘y%��?�;*��Eޖ�4N�ѱ�=�
)m ���K�߇�t)ߣ2K�������)�}Tߋ ���N�vX��$�	=�*Rt�MēEjl�#)];t���{�FM�lfr����
y������:p5E��!�r�s��y��	.mw9a>���������:L�{2}�ߊj���)�݅��A�p�k��c �ⶈ�,�m��Eٌm�]��a���Y�@���� `2�M�AD�A��$�km�G��c�lP�]ڇ�mH�����EL��,�_�n��,�Y# [(��c*8Wus�V	9?�wpX�28?o(�Uּ���)�)H#G�����7!<l�o֨v��m]���T+1d��*�ق;E?��I�2��}��ӽ
.˧�wsG�����0�m }�b�%����B�mf�ZF��`2�����y��G(��D�R� D>+[w��}2TA~���@�^xy�낤^�:�����=I�̷��`P�ے��$��W��1򴎂���/�[��P f� �ejpw�2޾�&��j��a�?vf�E�pZ#�#���/���{��I�g�;;��kZ8��?i#j�N���
�/' r����9ߑ�_G�Ҙ�Dܷ,�=4ͥ��J)�iZ�M��P,~�R��K�'���яh#��L�ʗ [�H4�ppWsЄ�����/U�O�ޕoi��?|��n$���Ÿa��вЀ�=��$��3�_�4v�j�����x�/~�Ԥ���_��+eD]e֤;�h�2A�'��p�m�� ���By3����I@���M�(|���p'��*�;�LUF6��tt1!J�^_9�f�}8/�C<X�&��������ì!"���6ܽ����Zn��
�OɹBE���r��$ٸ�V���L�f��$�>��'��_dB�w�_���Y溲�S���ښ����x�\��r�����c��O/�E'aFDa��"�c��ů�Cv�/�N�y.��;Cƌ�b���z��D=�����`y����;��n?TO��
�LW���^��>��=0<Z�s��O�F� �C��g�l�Zr�O�\�2��F����=�,�~
���/�;4��{�����GĹS�k�Y�K�*Z*��%0�m<�����2��߽�H)�������.�t��vk]�={h��.L���QU��x���%�������n��Z�2~Ԅgv6/d�t���Lϡ����'T�<Q���%}�gt������j2�����d�S��b5��9��*G!PKD�}&��M�!B(�7B#aډ�����bwj�+�!��8@x8�0I	-��v����0�[ha>)�1�_�Fr�10�6T�
�h4ؖ(���gI�Y!�g詘L� v��ڢL�e� P7!��c��.���~fo����2�2&�>�nl��(��iH��bs�O�s�em߅�r�
0uL�ܛ1������ae��%WW�h|���;�oHdⅫ�\��g��+PN{γ�@�!O>X|]�	��Ă��d�Pv�J�y���-��n�4Yzg����3(�7��bt�.�V,��pK�??����Ћɜt�O�k�!��5d�"T��M8���bD,'�p�[;�G3ǰ\�_�dV+jy���ɐǜ��ű&~��8�y�p��s�{%Y�u7$�����,K�X����_^M-����oǗ$��T��JW��q��fͺ��&D*�r����D�#{ =ϓG������Y�}X�,r���чk�zz]�`�&0JW�+��l���^{.
�lrW�"�G��u�� n6�fs>��T�߼�8����ݠA��d6����pzK���j2���g��{syqE�$��*�Ȃ���Tq�BE��>� R!1�=�q�B)�j� ��9B-�P	�	���Ҝ�<�ju�`��"fnoB��;N��a0�Mm�0x�:ME��Bɀv�ژ�\�� k���	u��k��PU����wh�Ϛ�ҥ�~|���D�X����}26W\M�/u�S�	s���g����DG��x�-�ٮ��8N���s�%<v�L�h!2�����@�RK]t�V�o}<i��9 k���f;.q���%�yo�O�K�#��t}ދ��\�A����N��E]��
��0�|6��4��˄-w��%������K�sX��0.W�W��M����#�ϠGЃ!�/J���\<c��J���Ņ������}�!�~��qGu�~L�B�I�
T*���L�W0W��@�=���z�*�ђ��jbۺ7�0�
n��~#X�6����ޱl1��b�>P���Wmټ�gK��7A9�`?��{U�&��� ��(;P�t]��s�_$o���Vr��T[lƽl5wqs�i����$C���O�+vٙ�h�-Z]�����b���$%]�0�N�kl뼟�f�A�Ax���}pdhC�W�	*I1^Y�LNT��2Q����5w�n�a*IƠ���Ȏϔ�ʄHt����۷h��=�lJx�!uO���UP�l5���x��R��B�V��#2!���o+	�������.���_`9�B]���]��ޏMm��������ch��ix��[*_��OO�{��@��MF	5��&�{��j2k;�k5�z�����Ṟ�9R'J��*	a5���uu1��ߦ��K�"�M������ '�)\<��j��g�}��)��-_w)�`cmO��&H���j�#��5�G�}���M�?�4�x�����_��c@ڨ��f^O���ƑC��E�J�����)a��eM��Wjشǁ�G�Q��F��c&ˎ���A���8���@�QE�p��m���1�s���"W��<����2lԛ6d��Qw1oa���)V$����l7Jc� ��	|ô���^�Q�a}�4�.�����˯��DevȽY�
ѯ��rO(A��.��(��im�k��[ɲ���Hm���_^FPO5�)3a�&D\ ����h���C�'�
48T监S1��z�W�1�{_^\/$���nd+E�D��@isC�7{3냒�����Jz��3(v��G��|�$���"�k��\�<�S�X���7�襽'b}�ڞA���O��h�S���z�|�ȇ��9ײ��_1�M���6kx��Q(��~���y��4�H��.F��m0^#ot%&�LSy���Jj�4�v�����>T��;�FX{m�K��T'#R�r��|��-&v��R�86S�
4��Bӣ�uJp�M��k¶�B:����G��_�D�ؠ��}.�%Y�$8�։u����+�2H(�|����@G1E�� #�0�f�xJw *(7!�f7���~�tV�T�	��'�>$��"7����
��������.L�6���u{#���P�qm���T���M�V�ə b���P�ކ\C	�T�Ǝ��K?g�~%.���O?�N&ڙBk4Mysz2ϪqR�g��7�T퍞�z4�)W�(Ϊ�,�(>�s3�P{�/DM������o}b�zGw�4J�}$0�a�ȧ���E�jux����"�k���_9��E�mڥ�qU��7␄�TN�n	I"���dd��%��	^s*�DTFc��%�!9����=ƍ�1�YK���"@��e(*h`K\aMτ�1�n��������\|@U�>m��+�Zϙ�|���q�Q�p��U�գ);TM�OJ�{�O�E��v�Px	~�
��-�����I�)E�ڋ�m���U
�ٵyΖե���}e�cP�r�C�u�Hʸ�����~�n�qR'�aL��豢�#DϏX��"ͲY��b�g�n�Э��K�R%�lJw����cS���ډ�#�#�~Z�el&ZC�p�G�]����^h���7k/�!
�V��X��%�>x_,�8�%����J�ݹ�L��H��[��$��f�j׀z��M�=^H�����7R�u�E͞�X�:�٧i8
n!���ݑ˖�i��e+}=���O]*v�g<�����*���� ���H�ƭ���@2=�r7A�1�3��O�	\����I#���	MBGx
�N�UjePӯQ̆!<5�4��U�g��V�13	R�8it�P(��񴻍T���|�}�8G0��G 7 ��۪�����.�̚h9XI�&�2Sf�J���+�;飶��b��o��N�
�>,���Fd;�A�a~6jL�������rt�����(��+P:�)s�9��Å#L��2(��5{Al����j ����t��6'�R-��s�8�EK/�fi���xY�s��MH��9;��LgB�:��2M�=��!4�9���NO�p�����N
`Hu!���1�q"x�����+BJ)�Fi�ܱ�ֲ|b[AG�i�4U�����}��]���3�v�=R>�x��v��*>���9�-)R��_y>�L��FI�LvO�VQ�e����y�̳[��i�iz(Zj�c����_�D��i?7�Џ�S��$�N�ҫ��\����De$ե�;7�� X�ĭ�pڢx~��Kf!�@��f�nkj�e��Q��<�'�c�%�Im�
���l\�����jsTS�7�5��_M��ՙ� V-#G��𦔟� �ث����w���]��R���^���ÑȮyE��1�s?^44qgx2�?��2S��1)RZ�G�$�6~��i5l�BD��`ֶ�OpGOq��(�I����tz�&���]X�s�+�X���L�f�xw~��o�IL�@�q\D��/��HG�P!�C�d[����IjAз_	K�˟�,��i4r�z��� f���r�h��v�"fe�O�n4D�K��M6��U�f0�x������ �ǰaݷjls#��+�ih���%�5�`Z�l�G-*�Nw�Q򋺄B�VrҀ��Q���#�I<ǄOov��C�\�~���.�{��S�HQ���-�! �%&��	�X�׭�ܭY`�͕^?r7�?LFQ3��VR]%�=���!n»�Wļ��rF)rB?1NR��L�� ��$1H��9�	��<�G\�����)��ki�D2�R���ԝ.F>0�������h���[U����˦��W^�!i��F�Y��% �RNEĭ��������~l�f��I��_�f`�($�|�%����d\W_ZF�+�8~k��x$<�4��D�짪
�x4�K���pW�t�t>D�2��a��� ����[���+_�ޣ�/a@��4!npgUp�Ä"�K>��#�s@������GW�����ϒy�zӦ��F���G��+}�b[�k)6ɗ����ZC��,me�}�$�o����"�(�?��tL�`�ؽ��y��]s�пƚ ^�~�өYJ:�ak�n�|�Mk�I��	Y�\�]$�a=ݟ�}
��qԙ�q�X	"I��6S{��V'2M�Dd�X� t;\��YҪBl����/Lߴ�m� �.߹�A��*���5��W�xP~%�H�����~2��J�W܆n��<%~��7�"�M̪u��p�X�"􈄅��Py������>\s�1�6�t"����1�د98j��S���5�aZ
k�QN�g3����[�T�%���E[��ڣD�S�{H��b���wC�Y�1��˼ӎ����S��ty�Hc�I	��L���f>D���F_��#��U5�� F�w��>�t��7�6_�-����lHf���1�Z=�+�lv�$.Q��[�<��a:��6ʠA�Y0e^{���Ŭ�J����򧙮���xZJ�"�r�L(´���������+�7*��e��&���b����r�d��.�笑�Ҏ����d-m,́ ���J}�ZV�%G��+|ciG������}T�x;^@̖H��@������L78�(0�K?(������2��z�<���d@���}���{!^/��݃�oZ��=��G��4҅��׽��`Ifq�;�<CZ�pk$Ч��t�]��{9c�?�?���X�%Xq2�(�$������I��K�CS�y��R��
���#,입�ʌz~�$J#pM�	�8X�A"*�+t`�U�/(nOeldd��
�7q�E�S���dAwL�Y��恣WQ]`��T#H��`��"(��`<�b�cᦛ���+_�,{���P~pߦ�;����bM�0��6�W�u|,P�&غlnZs�m�Dt���U��.���(;=��:;��J^�i��	7F
�,��}XM���+T+Xz��%��m�~�g�����E�1�^�.��b�aG�`}
�\ ^�V1�e�����,z��C��6$~`����X���������}"�gS)%M2��j��n[E(Փ�c�2��m��?N�p�F��oV�L���a��L1��l�N�ϧ��ʹ��͐�`���lw������t������9�i#[�P�BM�Ϝ��2��1*x��u�&�ᷔ��}M�Z��mJ��A(�:l�h
���E�F�D��z��U$-�3ę��Y�'�D�Eg���0�\x�昫�ۺW��B:{���%�e'���2�۔jӂ@^��޵��i',�̒l����ԋ]��#v׳�.�S,�Y6�hE�T�����k�P���ˮ���1��H����  �9g\���r9��,��FJ,'S�����R�l�Μ��H
w��^�#A���<{f��kX��q�#�5���FJ[D��X�>9�C+p��̢m�"�ZD?���"ω��Q�_[L.��eI��>�mDcȺ���;U���r�eȢ�r�*�3�@{�fެ���[�5f8}T�����6���G#
�����>a� �K>�����	b�f�F��J.�D�t�ď���)r�h9b���<�p����<�dP�A+�� �z�x���<G����/��1YM�f�ҩ>k�+� ���z��D 8@\U-6Ĝ]�B>GQF:�cås�pn���S%��1 %+!Е�WG`V��3�䚘.�8�z��6�$x��5�O��n�z�	�7�;�M�Qٺ���<ķ�or���6�k>���#�YĚQ��>;Ȋ����5֣1�Wftݴ�h���3���t1	�wY=-���J��?������E����T�<�l~�1�0���6~�.*�%U9MM����Pz��G������V�̿;�ң����\pB�~�����O��>�A�C�L�,b�i9I�����5!�8��/�ج�Ha�£M��f�.ߑ'mȾ���e��~,.�b��8T����՜B����C�yŴG���m[�:�X^�mѶ_'8�Ese+���g�<�G�"��M�}�&����¿��mMk䁖�Ë����1: _ۨ�wO*���b��ezy�	�>�U��.�T�CР�7�k��i/w6�9�9V
�E���G��r�8��|N�vn(��u� >yl
i=�U�i�s�,�̭�*�	\��c�7��EBM,�t�O����A$g��s*�yA��$���l��'�6�6mݸX�1��V����p}^t���3]��{!��9��ܾ�������&�if7�/�3eU3#P빲�M�8C\ra�,�dPr����/5���n�J!O�k
�\���#��ޒ���Ӈ�_�|�XV�x�n�:#�ɇ�As��'��av�_���'��f,���<�A��E��Sd�N����1��du�(�^�Y��H8�l_%T䭑�~U$�%��^��*��s7h���N���H���߮ٮ|M���+o�P?1�O��#�^&i�j  hl3�"�6���C���e4Ppz����Т:�(��)e��x�(��� t�=��GV�s�j����h�Ov��>������ w�&�����*g���'!�L�pGo��s ����,Jt�!	�lw�(K�L�vA���M��>�1d���O�cJ�&�/���$k�c��N�Mn�{�__盯@9����V'#�[5��l�J��Y��H�@���g�Q�)]
�`Րk֬Z[)|53j=P���D���ń}
F),���|Y�����\�@�f�����bO%;���n�J:lk�r��_9��%��/���u�Z��k�KC�7��s�V�bt_����j g���=S�q�ҹ��:��=��� �#]u�6�F�H�{ji�*�sR��0�2b������7��(Bj_$���G�'Ak�eg�f�g�҉���GS̳��8���}0�(��\z��ԷR4[�j��sB�8�)ua�hR�:+=���f�������1�NY)�{b�C������4�_�3�Ş�����F/k��*�<��owsW��_j��2�t��rB�̏�x'��z*�^��U���j�dc��&�^��:_Kv��!*�l],�yAP�\*�E��7��e�L��+��<��&�K��&$�����M%0=`�*l��t���oت̖ZV�C���O�H[������'dLm0�x�k��C�,����1X(����D�}�.oYݘ�]i�BT��ê9��l�Q���c�4��:�r	���ˏ��3v�<q �c�20̴0����dq�SԀ4�����ug��h�{��D��}f��Sƙ+��'�I,�T���^�1vv�Ǒ���7�4�H1�A-�~^U-�?���@��S_�s8�c�9�n���)�<�����'m�~�,Ԕ� )�&|U��Ni�7%��w�K����\X�!K�m��,z2�_�jZqf�2C���T`r�WA"Uk�jz8��y�}B'��i>U����UŌ'���=Ld�pՅ��q���,����\ �kx��QC���B�p�f�Z�3p�JTD���/�� ��_ř~�h���\~��c�������wZ��hK{�q_��,j�`��]�Kw!�ÿ�o���X���`/�,Œ>~v���Ixa�ϵ��� -�Dz��$�"�ܤ��έ�=������7b��%wc4�D7���ϳa{�K� ;*}n�MJJ?���>o�\�0^��T�-�c��+�/�9ƨ^3���ƭ�����tq2�S� ��%�W���w����h���,H��c�~��f@&5<0��|k[��d��W1�4�9��GH]Z��k�j�TgVf�lgz￷j�C%tH�^�E%p�e�r~���J�b/����ڀ�C��D����(��F��D��E��j�9�e� ��l�D_����� _d��AL�$|zǆ3f-3�o"c�u\K��B��2łJ�7�_H���:�,<7._Z5�(A���N�䵦�4��52k����yf>$���^�[���i�����b�x�Q�b?`K�knyR]
�M.�Q���R�8A�L���7�9S9g�M�W߁�>5�Tl|�����e�CM+w��c\b����H��L�%\{�]NVctpyP�������t��B�NU1�h@=��:jR5?SS3h/��oJѰ��z`M�b]���{;e���W��f��;�ɔ�VOg�r[�4�b䊈*��_��y�q
n�NԲ��
�[����k�~��2D�tƫ'��;3�G��Y<vW�v�@�S�A�7Y�{-��i�dt����i0G�� ���4�N����nB�~�;w�nxn�"��KMFv�$��O&坶Oנ�J@�:=������`N��Jk����х$��I��H<{e[Af�����P�8bf��Y��n���`Gg꽱��R]9�9����˶䮂\�+k�&�U��~���1A @�I[���RY���d���m`�-_b-�Qom�	%���y�-���B�^�x��L@���Xa�Oz$+Ys�yn	5�	�}����J��h�H|�\�S��Q6˥.��U�N�Ood���F��{Z���G�-'w�ٕ���n�Θ~t6��R��k}�������'d��A�րP����*�	�'�z��o,�n�8Xqzx�w�kg�����9���<Ape��ݘ��I%��i3L/H�ǡc���;��!�l�U�M��Rwą���g�>�	�ڜ_�F�1}�X��d��YJdaU����gO�_W�]��`��m:�"焻��L^�k�|6�^J���" 5�%I�r�HZ���a׌BQ��[���T��>���$�����Z�-���F��
�P{�E�W��P�̥B�I��Q���'Ĕ��&�tO�0�9��S)?U7*�!��g��x3��i���0����홛�l�?a�;�~i�����jUU02�W�Z��V[�-�7��EY��į�{��Q����q�5�~o��\՟(ú�S�*F�o1_^���z�;��к����tM����7@+;�-��oi���y�N��ي_h�9v�������(�arf���!�SRI����04j�K�R>~ND�kÈ�ƧtZX�E3V|�4�5z2��f��z�K�!�'���-㖻h����8��vO+>�N�0�u�E/һ=�ʇ2j�i��f�1� v��4W=���'k���/p5*A�e�w�ߐl� �]�
['��VJ�.��y���/g�I��нt�t�s��2j�!t�#�;X�an�F���vb��o-��U�"��[�T���G��c|�W��3�_����y�A,	��zΏ�5LF�5_�Jʀ��HL��z��wI�����Y�r�":��,��A�q�>iZ$�?rڻ��b�Os�������Oc@���>[_��z��ݲKa�8�1��bs�6�f.��4���6έ�G���!��XaA�|��r���na�l����rUI�� ���H؛W�A���u�B�Cn�/�Q�QD��x
�n ����A�j�<O�3llxb��� �	#h,Mt��m(8��o�F���sj�=�'�Q�/D_�T!��@n�%o���T.�pY?FC�M����Ԓ��vJ4�Y@Bz�~<��D9Wf�IE�
�bt�>A�
C����CA���U��*��V`��	W�ox��j��ƴ/J��:c?��d�����;�����;]EE���.M��Q�}���u��J��,ɴM�� Ѽ�������M��z�4����Ȥ�iO�|��²�P|R+����H�'Eh;�ǲ~F���v
YTƩ�I��`����|��h���q��o��o:��;��Q�$1~����4�� ߋ�A���Rp�;�`���'s��h�"*tZ�3)��'��3g��7�+d�,���������"�:��m�~5���Q�\��SK׊�p�Z��ذ?:HI�X=���K�ƴ���}_&G�ǲ�n���m�=���J�IM4���q�E+$'�ʦu�H���]�B6�(G_�נ���y�)m�������$�g�?�(C��N%o�ٮ��V5?f1��6�y���pqn|��B�������>�a����V&�q��w��+����6�;s��îS����/���?���4�R�������*��"���J���>���P�7���)+�)�[���+�is����EYD6& ��E���t����7�/���;�L36�����K���G����9�%¡���]������4s�h`�v��q&\�\�F=j_��V��G,!z!�_6]�$CJq�Z���U�������{~ӭ����,>�bGe,��3u�` ��kή� G��"`�c�"�	�ٷ��)h�L�0�v`v??O����l{�V���z�U�>T1
<�4�6C'�y��>�Q�-�uAπ�t;���U�^�RHd[�f��_���4Z8KO��W��8�>F�h�a�&`u�?����B���<6B��%nnj����ը��`��d����a�2����,��'�dEF�?"�����-k5�^P�)Y���P)�_�;�^��� 7�~6��tG-�m��(�δ����̯�[����A˯@�A#@�v��#�7��t���b�����^�C�
��A�	��W�3����D�J�#qd� $�n�\L�l��E�%dM��j��&zI~�,���ퟁ&�U.�������cI�Bc"Ҧ(�m�^��~x�:�{i�V8�yI�2�{��Bт������P��y�I8{�X�BO�h��h���yEa�ۆp���8��f���Y؈?[�0�s�(�K��L,�Z���R�(��Mj�W8"T&��5l�u?f��g7�v�r����#��S�3��ޱd�o�Ve��`���)��~��;��m,�Q��yx����K�.@�`��v�]N�Z�1�n�5T�m;D��4��<�Y�(�A_!����x�?5����,i,j���Q@v�@�D�Y�O���j�h�{5oԆH0�3^iz�ލ���`0䔾��+7.��u����5�P�T"M�����T_��1J�3ˠ]�	'��cl��������y���gm�M��c`XGK�w���c��0�R�"�!`i&�uC����,xXsz�p�B$]��� On��*<��MZ��j��W��`>�K���� m6-����[��ج�����X?c:ea��9j\Y���7�ul��;X@d/�|�0̗h�c!xq*4���CG�ۡU� �}g����!BM�EL�9���
:@�H�ͫ\s��m.�u�Ƹn�f�W����/�(��	�r�q�㴜k.e��ՀkũIr{ٸb^��)s�|OK}=Юv����3Lh �u�l�jV;M$��Oزu������D�vbY.���Gľ�%8N���աg�SJ��gM�2���k�6b��o�ӭ���<CXC�Ğ96'L�gF��*_�/@�v�;"��r��V?Kfj
���� Q��F&��2#����
�ty(�o#���ؿ[Q%���GR|��W�ڱ�N���)��~K��ԗ�7;�B����S���Ai��YD��F	:��-AM��5̟�kiH��I�m/�M��V�`KYsW�D�۱�6�h$^�?���s���7	M��#�x}� ���ܸ����u�)�\����\�%��t,+W�K��D�^c[$�kId��󁂆Do���W&g.��W�S���dO&�;�*x�)�����~%����8���J�X�Xf��7Q��WR�ERa˾�4�F- %�k�^���2��@kF[q3LQ���t�1U9��K��nƘ�����E�<AD:��W"����'��&=}��&w�]�Mt�T�:��qZ?���o�%��]@PN^hE7G��}
d�I��`~A���C�2��A��}״<���a&������i���=*�6�q\�í��	ӂO�A�!ܪֺ�m5|�бm�ŰZ�r�b��k�A�vE�O^s_q�QF@�Fd��y�ƞZ�DY,B��-8��}D�j�(���u����lQǯ�Y�A��+�ѐy�^��1��]U�H�(�Tc��S��^�F��սw�AA��1�AXF��"IG��H�Է��i��vR�o�4F��_QAE 6�|�z�n��N�V>kī��9f������:U�cz��k���
P{�`鲞�Tf\�X����{b
���kqK�4	L���n��M��i��W7��댊���>�WdLw^(��(b��PO�!�������h|�s����������K��l>�޷+����30im�?�se�(���x���y{�Eņ��<�x�+�Ln�~Z�j��|c��%�p"Q-�Fͽ-��:P��H���Ơ�C*��ag*�f{�1CT!�C�gX�ؿc�']:���s����L��ő8e��h����ḏ<�D!�n�I�Ґ�6:�/��"�"�b`��%A����4L�� ���1G'\�/��m
�+�=k%�� �ٮ�N(����5%@�X�7�:�Al������bf�'; �,r5N��
A�wE�q����-�c�k���ޒBiJ�򺲌�C�ZB��|p��꣒��]�w��(GByr�ѐ.!��M���4�WK��@n�E�Ҩ��/w�,Q�[	��N��F��/p$i~��⹍�J5���4Ȕ���z6����+਎�꡻V���X����+�X�$��Z5�;>I�-�����S�9.��߻�_O��ᢥ��W����|�x����\�M65J��}��Qo�W56*!�����5�I�������R�~�u!F�e�҈4;Ρ+\�t�'����33�|㕂7�[�x�˲�E��0U�|-��E_%w-MZ�o$���p��e�0�f�/��#\	MCO�������Ah��Rs�e[�u��:Rbw���Ӂ�̋��8�0��Й��w
f�YM�F����}ݬ���r"P�私 Xo�}�	�X�`�.�5g��X̫P	�W(5_ݪ�t�Thɱ#�%2�~;��Ʌ !ǣ��x��]��ҝ
�*����vF�����y!^��_NA�����k�	�}	2�M+[5e�*��lM�۠j�QSR��
|?�� Om�K��Hw�I��
�^��Ԇ�� ش�C��2&�Zz��Pjq��H`ٷFl	=����]V�лWu$`-G�*��qρ0��(��d�����/���)�I�?�ܣ.�� �-K%/���p�@�w�פ�Z$z�Y�c*�^$�Q�~�D�"%�u"^0<[O�8�>�_AYj�ЫAqv�57 �q�hS�fw�}�X|��2��V�u���ov@d���Cӑ�Cu�Gh~��C�<���T���5Xb�2���#!�9�_0IFc���tR�ki��N�|7%6�/�����]H}p�*癒6�����[���{<���R �:��P��ă֍�(�����hѻ_��H��=W�(x���r��j{/��]He�g��u�Vw�r��` �x��(�k�+*�݉.�/�=k�t�
����Х���.�j�U*M�ʰh�<;d�k�9z�<HC[��O~���k
��۩�(Y�>Ioo\����P�x�n)9R���Pԗ����ao�,�_��j1y:���2bN�`�>k�`�-�C�ovw�s��P�w�AW:]�����`�Q�ֱ��c��_q����@A��_��W��9(���E��������t�J����5� "�&_�M�F}��~���S�	\�(LMgw�g�F�
0��wPi�.h��fkۜ��+�K	G�����7�Q;(�ꖖ����U�#���ҩ�(C&=<�����8�z(���!o�Av�L������o����9�7V!pr��~��r�JRs�T��ۍ8n��V�}��Qb>-��(�,\�*�ܔX�#�
!�G����fj�7&l5� ��m���}��}�5��6�|(�\l�U��Ɂ�2�|Q�d����� ��T�)��`�'��fl��\ܥ��)�M^.��k0L,�{%>��Ә������]�}��X��i�!Zÿy�eo��9�S5�e R��a�,{�������2�/+�w�R�o�f�d8-�����yl��EN�B0x�OvH�ͳ9Q�
��"]��JO|�##��S�D�D�l�����I?�����O�C�?t���8�@C!	�=q�Vx܍�\�Gq��A�.k ��+��>�f�������*͉��Y��o`�'�<�p�T'�1��J͠T�&�/v kQ��i-���,���<t�eS��x&Y,��vض|[�
�@O=�v�Ñ�S�Vt�'}���"М�(�2��Y�n~�3H
��>Eɂ[��,�ϫ|2_��F�T뗕b��z/ܨ�"K���$�r��p�s�H���Tì*Je�m�I�be/�m���<��R�+"��ۦ�b�����vqD�g�#��/� ��0�^+��1S\�&MEϣj1W�K;�Ai�����üL�n����h� \��X�(@�6�ڑ�I�F+du��ű�u"'�@>y� �ު2��,� ��~��R���3��={x�^�U�1#���o��]<�-�R�LI���*�NJ�'U龷��j��@ػIl�w�m��[�c:�n�ۿ`�,VOL~bR�д��Y��s������[S��G��.������Z��ϥ��C&Xg-��
�R�_q`6�IER.O	>B�-��RD�N�w�@~ ��ŭp�&��)�7���u	Gn��j��7ԬU��]�]C��=�i�YWz�k�E�y
Z��&�#��Az�g��i��r���9S��}L��3��3ު�+(�3�❡����6�] ��9��L%���s�#a���'6}�s�SV-��E�g/�C���b?���7a9���#L\���<�q�n��"��ѳ,����YJ���().n^�C�!��A!�+F�o�:��u�|���J��)i��Jo2�ueh8�(���H�yȖw7����Ѣ��B�{�����~>T�5T�.��y�)�#ǐY�N���a����H"=j���SQ�o�u�S�ʚ2�av�4iǁ�z1��ŝ�g����9q_�P3t�hn���Yr

�96)Q������h��O7�IecO�k1�I�%���H�L�Cy�-�6EɮҪl��B�V�ֶ1�9ISS�FFJH!��=�����:p�����������r���L��C%�c�����뀊(�ӭ��Pe�S�eq�L����?�JdRT���n�V��*IBa���&s�1i��S��1q<y��������@u7ܶf����Դ���SB���.= �A�v�oY����ʚp��>��%���6Q���;�������"�2�O�m\�8씣( r2MLF�C�o�7��r�Ic�G��"ZuZn#֡�pl��*ӯ���!��-]'����1;�Q]�*l]���h
3Q��|9<mDr�����.�d��,,�x�O=�*�ό��e�G���{ḿ���w�1?��fMZ��\�}bn�X%�� ���t$fheߒ8����a�w�*:��?1�<>\~�=���N࠵r�h�����o %WNa�5;aIY��\�'\}�h\f`J׭�iK�%v�~a�?�F�BͿ��P�<X'�Ko�	"o�oG��Ջ����߆Ȉy8Zk��kD49���C>ŀɝ��Pw�y|m��b���`*|�^�A�|ߛ,����{���Sؕ5��:ú0��|	|�"���z�k�Cj��{�����.��&� ��a�U7��,�oz�#�4
������]�4W�_$߈�&��E��W�gT���@9 �T�BxT���
��Ӄ[%�d=;�S�k� FU\I��c��t��y��طa;�/��1e�M�n��P���0�j�ą��u���ٸ�&�����
f���:�mF��������P(a����,U8^�؝������F��\ͼaa�`�lL�0�&4�'�eٲp�ήqv#���?���5�͓C'.���-��8��3�ɨDjydO���y���I�rP,����7N�oFv��P�ˊPq�	1�g&0��gl;u������ h.p�z�������K^�!|W�Z�m�+�6Ck�/N�C^�Т��v����5;&����^���ݦ��*,����;�?�Ӧ�J��.]C_It��\r�`�y>�ըb>���.��p������a���4�A?R�)/-,��53�:BF6"����w�|6�|&fc2?�U=���Y��K�8�JU��R�yZ�!�I��lO�^��-u�I�
r�Ѿ-�9PD��P�#�\%��n�C�͝��s�7|�'/���+���jr���nr��L�T�1x"���T	�M�w2�j-�?���疵+v`�ib$�e���w��r����������T�uܘ-ϵ�+��Xt�vn'�ԂG��0�q�̾�V��]Eܷ����Q\M������pg7����ߩ�/����[2�1�2<���Y8����~�} ���H���N���Dxw�������{K�Jk�m;t�3q�\��CK�U���u��:�C#�_�y�S�D��COn)��1���'��N؃���<D+�Ksș-�����ui:��``a�l�H3v\J���jH�G�+-�UϦy>�_��1���κ�Jӕ(� 	s�m7��;K���a��dE��1l�~�Au�9G�<~�7WpY�3ҥ����Ij�4�nw�ؿ(�pr:kK��`T���
�c�ڤ&l���C<�\����d�af:��+tL$�ƈ_\?X����E>l��_ܮ�x��ǠN���E��&�JbR$E�����Y;�W�;�v6�
�.����^D����j<�<���pbo��h�������}܇l�D���)��5�֗�
����/?�ſ��[��T��-���F�4�����7���:�b��@����k^�A��t� �vyXב�{gg�>�ل.d�e����~?�u�����$�g%��/��y�^3�����,�z��01�3MRN�0�,��r�2���a󸌠r��6/	�O�m�٣�C�W��� ��I�LI���+����)%
�de"�Pb�$i*\ӵ�p��9������(HǮTO8�@�NH�~r�+��$�y��U��*�O�jq����������`)%b�o͙�bƆ��ߙ zz��|�s��gL�$��<bˆ�șC�I"o��xĊP�</#�!�ǚNf������,�u-�w �-�:)�_Jk�����uW6{��]p�c,�>�F�a����m܄W�k��!Y���G�7!}Q PU4�>���8�Uw;zq��d�j�V�I[ЬΡ]�~~�C\�4��c^�疷8������QѼ�&t���P^~� R�֚S#�"�즖��m�=��6Cឍ��hy�.�(��0i)id��t.������Q>K��g�IC�M.��۬K3U��;/��H��<�^��۾}�~�3�{�ӯ�z��l���.b��ol���Tj�=�)K��TON�VP�n�(�����}�R�ֳ�|�����S�[]m��iM{���Q���yi�+�P��Y^���_����O���w��R�ZTMm7���\������̤3ɏR�i~���E�C��C������i����
�
��(Bx�L����Q{C�����B2���M(Q�";���M&��86,i��~-M��G�_�A�WW���������*�6�Λ9f����Ǫ`���Q_[�/�%0Y�����sa)v��]��1׏��	�?�1'ۢ�c��D�,�*�]4���'�
0Xo�1ؑ6����E�a�� ;��U���g'@Ogbu�}V���&�j�5���%��䑱�"�dfD�V�����n�,bIu�_,գ�{�����ܳ�v�w*��t�̋���1�l@�
|Z�D/\fth�y1��l��jG��3D�#J�U�x������RèyBzG�n�!>��쯮�{�\~6_�A)�ƅFV�d��;����4�%�w�R~����U)�C1_��
���g���Kɒ�Y��c5s��[�EN�
���!�y��ͤ�Y`��aDk"<	�3X؀����s�|�]������I�QL�Q�m2¥�����y����?��V]nA��Xށ�"�Q�dv�H�FH(.��fc��s
^�:�a���	���ݽ������ ��밟�JaԸ��KR�I�S�0 �H��k�0�kK�|0<4�R|�����=W>Sh��]CX0��8�?�ϋ�����1��E~ޗXຽ�i����M����ّ�֔����*�	OAE��f&����~ګ�q���jR"X��Ґ�C��� ߨȑŴ�K���}��RC���,�����C�W��hF*e�,���B�Ԁ��
B�D��6��j������@̍�M�_�b�����>�^�H����D���,|��G��͠�F�m�灩(r�V�j-&|�֙V�~��GB����UyY&�'#(��u��v�T`}�wl����z��m�j��}��l�}�\�����z�
2[�3p�y9�P"?ǜC�.����a�p�<Q+��(�N�Y�c����v���gVᢳ�DJ�E�CJ����y��0�^��7��è�|j�Hȴ�A������Bg����h5}%j�F��>���0�\d�^�ȁ�����$�\2��+��)q}.����w<��]d��>�rt$�c�f�@���d�[C8��{��|�Í��0�T��Q&��P%�����d]܋�_�zٖRm����k��׶�ao����pE}3�&J�� Bڵ�J��֒�gEd�X��J	�y����wnw	�7��"'�;$#L��ٗ.��v�SS�ய9+��׺BN�����=vb�_��ҫd�x�K�����ݶ7p:?�}�`�U;|����ٚaݴ+r�;�0܎�ÌR�v�x�qV�Rد	r�D���� =���_��
�8���]b��ξ<��ϐOl҉�?�!���	�	��q��4Je��[-&ftb�w�y"�=��3B?]�	.�����ׂl"�����Y�>l�A���� ��ì/B|؃wL��N�%[YY�	�{��"t^O��/W>�dұe��+���A�T�S�C��M�G$�R"v�a���3q<�~��������F�(�&'4�g��-�Q�[y�>�E���&P�Z�V�ӉU�ݟoeRAi�\.��J�SY�@��ϡ�K��|��g���&�l�)�ŋ�"�������������m쉋�!68i�gPwߢ}\��%a� g�u�p���|JlS�{N��b(�ʻ ��sA���n���
D����2-�����]$����m�Y���jD��Z�E�
���2Q@�h�j������"�䇄9!����v��[%��~�%�V�ZA'G�o�yMy�^a����;��/���xg='0�Ȇ�G(mAK�R�K�~7�=�ۗ(��l=ձ-�2�m9����ǩ������H�a��{Xr��x��*��`多����iJ2���R/��s$a˞�����W�f���	���N�78m ��U�";����9�R'
W����eC���0�Kb�i-W��I5tHd��
 ��/���6E�<R�������&Lk�3�6w9y�1U)|���E�؊'u;���� �W����;NW@M�����.�Z���Z�pu�4���9�r9� D ��]ԃ��9��Û���xHl�p:�K���tB��'�1�B�9�L�[T��7k�\���X���&��B%�<��������aS��X=,՜`��6�?�6"�	���ę)�R/Jׄ3(ki$�&�� y��1�7��{�r��)��pd���}�I96�kl�@&P�l4���7B��2;�����ޓ����0�3�m�F@�C��}� �j���Cz]Yt��$W�2�{w�7 �>��=��P~]��2�� ��S��7���Y{��r��/�!���Z�])K&���k���[�5�<�7��e�'� Rt����4�='e^��KMw�Rح;%�g3���\�f� �`� ,�j�ŭ�!K��wJ�����\=tr���'��#yu�/	C�3&�{�GZ�Eٙ��<㽑�ݑ��1_��+n"d�*R���]"+(2|,mb֒ꁞɞ;��ܨC�mz/{�A����CM����t�nP ��r�@��쟍����^�LM=�&�J	(�hA���6�]D��1�� ���t� �H�p�9/�kfk���J3���-օLQG���D���k��@�6��b
�ߺ0�▋�"Oo(��!ҧy0�ֿ"|�����+kj�6;�Ba��c��a^Æ5?����������N�q���\�!�	Ii��a�����rl}5\o7����!�޲˫�K��J\ ��
��c�DQEla��?
uk3μ5�;#([�]�f����_���{_]���Fv�� xj4�3���S�ǂ`��{7�pj���8� �MH�6�,�Io78t��Ӏlc���Bv�X�����P�@un'e��q�-�	ܲ��䳭� x>�4�s�sE�TSb����1�]��0�� J��M�3Cf?V$�x�q)�,B�h}��,��lcy�2��M2�ݭ�Ǵ�tH{ַ�RȺ"Ѡ���O��z١�s���"�=���๭��Ռ�
>�c��Nl���_3:7?��U�<���}��G<}T��_��&�����3�R������Q�ΐs�m���T��"�[L�	��G�CG��[��kN1R1�e�@*��,�i�s���0-󸺰�D?��q6�.n�P[���$����gnE�<�a O;_P̊<f&�>U�a� TLR �� �ut�|�% �A)��E����ή/լ�bƸ�J��r7�;���+:�=�~��;���cQ�gb��ы���D1t�
(/����/��i
ah��B��+���<���@��bƍ�ؒ6$�W�-�Pk� ���"U|�1M�����ke��{8,|�;�}ʃZb_<�@#!0��' ��@���U��r:'�r(aX,X��U�z�V�(HN�I�h����|V� =Vk���Em}���5��k�l���"�i�c8�ϺN����
��Dʌ̶쎽����H��a:�J�A�#V=�����L/�{�Sx�r2[/r�ʹdRH�An�k)^���C'8��Q@�+J=�,g/�*y�m�Nj��b�T�]��O��A�h�bѪ����尠ٳ�� ���KevM �,����<��)����|��i�S��|���V'�ԝH�n�-��b��얙��o����q��/8K[�d�t��)����HA3�`��@�K]K�T���E���ʭ�+���m�&�켟���EP<��Π��O���\#�ծa�[:����>��f�͹��,n��̬f�����d�mJ�%е/dZ#�)����0�{�x��lGr^�#�,�� ���	m?�:i��`0MX!5�wq�x�2K +�-$$�WY�Lp�ǧ�P�2���Ɇ�?�W$ׅ��v�����M�B�3������1�ZR`8�Wg>��l��ȍKJ9AlB�%8��*JB�6�/��!e۞f�A}Q,�$�X����9'�l��l
�V�ȴ��kY����?�26���͈e�sw���~���D#���WC�o�.�o��7�~�d+��0e�*Bܳ�.�X���O>s�{(�a7�=�[������3E)O�Z<��aS�ܰ�ڋ[L7+^�ڡ���}q��y�"��]G�k@[�15��]$��0�ÑE	��*�����8��)�����=oުɮv�qb! `}�Y��y9I@�,U�"iS.�
P�� �/to���ﯟ�bd��&R�!膕�[/��=��ߚ>�2�����#���]�v��ɼ�s�y�Hc��"l!ˮq�4S�6Ϛ]`���y�����;�����+vX��
��1y��#Y�GW���B*}��|"0,��N<0�y'�&}�v���t�g�M�����w��_��#(��Z]K9���j�-k�4��83Z׏F{�����z#�H�A�D�r��������C!�ɔA@�Kl��s���2�p#Y+\��Vr\�_�w������R�w�h+�H����UN�̥�6v���WZ���)�+/S'���|/�x�jI`E��R|d!V�%��;�)~�9����?*����w�,<������P`���0�թ|@��!�  ��`a9)ID�q�S��_!C�,E���t�tKW5�y2���҂:�h���p�h�uP�O(B��|K�Ldo+MZ��"��C����v�L���u���:vR���j]�V��-�=Ah�Q�V1�s�Z}7�o����2���aT�x��jC�$Ү����q@��\���Z
ZO�ز|��KW#dz��4_����>f��nK}��y2G������#��^i��WJ��1J����o�"� �ªΉ��l�����?��&�t@����+-��Y���+c�f�n��W.㖧�]��w�g����j�Z9�ס��y��k^���]2���Cj���&�t�j-��9?��H�Bk��Xl���Q|2��!��0�4q��6���������k|�Ny%�'�[��δ ���~����wPC��M�P]P�U-w=�4q3�H٘{	xзpZAN���jJ�a_��c��H�H;q�񁓛�bY��J�j����*"�(l N��C����l5��a{h��d�4�k���Ć� �Wqh(�H��ZŨ���6X�Y�W�=b��*N��{���c�� �^�~�Tg�z�2�t��wǂSݘ���?9Mro�D�^�+[�>�ɸrr,���j�k9.)����YK�W���e�*㾭���g���Ԁҗ��u�wW
1�m������ĩCb�46�^��h�Wj��"�T�6o��!�T>\Y��O���.gb��6�*�0�?����,�SYMD�:C��bޫH���O~~a}8�e*�M8l5��Dh��\�4���X1aԮ8be!ޥݿ�4X�򿱾��^�Z����9�c=&��o�81��ߏ 9���:v�z�0̮fbe��-�9��V ~���ܜ�?���CE"��a���k�G����T���b
(��"~�����-��	��ח�"f����#;��5��{OE�(#6V��Wm��� ���lB��A�f�cW�Z/�p�p�y�z@�4�*���@��.�p�d���`ڴ��&��;v�$C�-y�)��]���y�]C=��$W*��0u&��m�V��0�R(��)�no��|���]tr�Z�NY�%�#J��2O�����h~���9��'*���pɦ�q;�(���vQ�|J��QC�zx���E��8��}�Z�o|9�� ��� 5�t{��~���?[��*�k쿏T���T�GH�#<�;fe��x�v�QE7�k&l)�-a'�ydak��*��N�V����d�P�ӶP3y�ΐ�Z������gauo���,1������h5��&f`(w�e�+��h�=�1=;;�����9=��E�ͮFhΈ��[�P/�BHd��!���:����^Lњ�������Ax-��d�1UK���� i�ʰ9�L�?�l_X�IӚ;%A ���?���'􂯟<��]_�C~��������t�5_�N��xK�hF���^�`�jø�,;�����������tGƷ��
?�VJ������������'M6\����� T�q�иO��J�p�9�ĉWɹ'��F�*G��E��.q�"�H�n���4��	n��%g�Ak,=Y���	o��T�c��z<o�E?t�k�R}�9��/��w�ɽw�o㠻�S�kd ��,k�al&�q�R����>�S�йN��RG��lˣm���ߺٵ��vjy��	�aK�g�ݫ�C�3��BV���}]LC~ld��1peQ[�$�jq�t@��h=Ɓ~�kU�<�H)�nO���#�b`W��$�<�6dP�|J=��o�=��`�� ���B/n�)��.��B3�͛o���>�ʘ�]��>�0��Gk}oP_5G��mt���\t���T��4s�u��Ӽ4td��g*�Y��~��j{k�=��XP�ʬ'�d����ST�H�3���0c�O�6x�	W�1)�k��K�j7o�.'��+���V�{�B^k��S"k��둬��e!&�Վ�2���H�:�"�>����}�̋�]���<�v�a�Ǚ>�x�*����
��-���a'���������L��p���d)�.��^H�3<|c��~#'��jV�U	���lA��):B��-p���	s�!K��������M���������{����w�`U(X�&-���h��T4���~cF`�2��)����E������ ��u+�g�&��nn��2�g6[��w���w�s5��栓��֐�6����x�K'�0�Bw����	�NPI>�8r!0��}�W%�*��	��ۜ�gȗ�"�C��.�u&�8#,��c�x���g7�d�}�GԴą�U`'��ꇌ�iTC:���0��z�m} �ڂ| ��J��~S-�%;Ǻ�x�o
����㣖d�	���@(!9�12/���7�+���6������		�/-�[��wQ\v.�U[��:U o�;]�/��W�a���[߆c��5m�O�Acp"��:pv��I8��_#������.�!o����>�7P�ŧJ�����4#Ǉ60�o�\|&�hH�2��x�X������(v��Z�`@WJ�O��ٙ��!;Ƈ0�4�WԬC� ���Txx�=Yrm�PлuX��~�n#�3�`ݹe��6I��zv���7�^��d���D�m��R��2�����Pi�ޞ��cn�l(��İ�ϥ��B�2����<SӴƇt��vZ"[�l�o� ֻz���As_w�D�(��Q���>,��w||�	�s��|� �>�9��C�������5�IG�ϟka8mACC.����W�=(:Ų�9��*�������41���Q���̳C��+T����g�ͫF��ysP�<w��:�0��lh�n$
^E*�������>ⷅ�t��א��w����m��@�r`��+3����m��PנQ�����0C �iC�[�Q�b��z�no��r��}�^w�8'ȉ���sӷ=�`��3u�C�I~h�Ƴ4�YQ��l��-���mU捬a�O;�lo}�NSǵĕچ[lm#!�ɝ9cb�<���	0��B�5���6�w���"e�����&��Q4f*�դ%0�M�`,]�#G�$ �w	����H;�NӃt��g"�Ҹ���I-��l������T��^�!��kt���t=И����-���u�=6��n���\;�+B�Jl�Q_C!�P8�`7��= hAb�;0�J[q����S��*V��8 �f�~�9�)�>ϐ%��l�F�Em�+��}C��G .����O�t#�Q ����$���6���4Z��nqYU�8/��ӡS�C7��k�Z�ed��Z�6=�H�G�����C�����w����p��>I^�^u)���p��73�Q�kk���c������F�8��n����q����Yo�ӧSʻ��T��H���
V
(9u�Vt�T�;�qal�٩;B�^�����@F�#R�p��@�GS�k��9ja���-7��n���E����5���3-��F���؍-B��$�녌9��x�/9��$���IW�z^p��Ƽ��?��=A�mO��|��pȺ��wP�˖���0�n圃AbB�4e�0���/�����&���t��oA�E
Uk�@�'2\�3��gJc�)2P����QB���7Wˍ�Y��Ҡj�N����=ܝ��u� �BI��������߱j,�E䍬��d�M�,���|R"F���k�!�Hz��o̲�Z��#;����E���'����AS���Q!t�~nCb���w�?�onՎ�p�S�Ot�ڰ\B׊�X��hW��vGYeh}]YG��y���V�(����mK�C"����-H�á�B� 3y��h(���:k'�]�d���*��Y$�2,�B�!���ޞT�������|ۭ3���[*�>!�5yK �=[�_p�v�0�֥XmQ���]�b�%]�1kR���MhQ���u�c�$�
\j�eN>�;��u%Lf�QWR�Җg����!uU�8<��dD�F�7�p�w�W$�z	��d0��}H����_@�t���5�х�_Z��iv�F
��?��p��m�}��0�&trh5҈|�:Ê:8B����g��IwkB9=����E���P�K5'i�W��n���<Z�\��DU���Y�j.[a�Zg�S�4<�X��611R~���>ʺ��y�
���.x�v��W��8�](Z�z���M�-*�\�1���/���T|-�m���iB��]>p-�2|�5]/5f�:抛w�����9V�'_o�I�#jǯI�+)�I��2��?�w�F�_9���t����U�m��1B��n�kLR�{Rҳ�q8���U��K��QoK�wf6�`nzD��s�CB�����Y��o늂��+�X����c�:�?/D7�3���Z�~Ex�oNa|#�Л��>5Un��1���ɦ�(��y����5�⚤���@ �uMJ��PAJ7��	k�Մ+qxq��	�t��;;ܖO'���y`�C0s�^d�nzTx#���v���v���¯M���R��E�M�ai�XqA:q����A��MO�ѥZH�y���q��b��46����<��
�,�kNK�G�@�xA�H6��P��T��I��rAǃ��q�N��܎�f�
�O�]�m-uB�j�l�E��IE�7:���x���q��	rs���H{+"����ho�7���El�?�⣟�L�H�'��;���f#^%a��y��0��ci>DC�4�Y����;�F�Q ���֓w�@�m��X��[����w�]{�����.2�ny��X�c�3ShEQq��ݘ�8 ʹɐ�����T�#�{�J[�ȥnYG�03�A�K ��}��`��I�:-���vW�v��`];����ԈM�>���	Щ�n�ow��ǡ���t^2�ѕa�u�o.��\����M�,��K�H|�֤-3ΈL9�#Q��%
�YE4���������L�T�i�Ͱ��&T���M���A~���?甏7��[�!���$�Ug�(oFsg�����*��zEIM��eG�6E������[g�� XƩ�e��l�V]��^)D�c�0Wsz)j~tԻI�����?CH㲍�����yG3����P��С���r~a�).4��I:�Q�S�:-M���C'Cס�pQ;߹+]T�E�xxL�)+�M0��y�Bd�@�\}���yU��57��~%�_��*�H��][)}��rR�f3<��狀�=a�Ѿv���?��eB�4�(s���o6*�^������b|*E��us;6�XY�h�p�D���.=�y�����G����%A<���m<�n���h9KU��:F�pΥ�9v�VOn�?x֌L�@��A!�����u�)��xV�X��pzѠQZ�]2��h��f۞8�Z���N���Uf���h��� �%;��+�S[�Z���9�aw��7af��+��k�3��L��������:���!clbp�P)�UXO��<�����ރ��l[}��-: ����V�{�6�ʨ�wa��ʿEghYWىn��*�h�})3EA=#n��+Ŋ��u8���u���FT@�?u_��$���� �U\�����L:]M�q��<�tW{]�p�*�~%ޞQ�ʛ������ҒX��%B.?�+���o���h�\�j�^xe {m��T�,�4���~�0$�U'#7�w��lf�3��kSK��c�6-x�O�A�K���'�f�v:ݻG�K��%�K�SYECƥ��4poJ�#�xޡ��+�U&����������o>���˖B��_�](�����&�	�{��)#���'���������:V=�V�!�r'�c��	b�~9�_A�YAN��Ew��xh����5 s�����(ӄ���ɉ�:1��_0�=L�_0@�in����ۂ�p$9�R��i�ߍ��e������5XjDi���dQ��x�bA��w�
�V��^+�:�F���P�+#Q��}��lL�yFm��L�u7�OaX����K�g���h��/Qrl�i�*=������RV��Gjp��E��,�X<֧�Ǐ�O�K_��`����j_e��Nٲ��>�b#�S}��7a��?ꋮY�������[j�췪
0FD4��޿"N�a��N���g�
��/��șOC[>��fg'fT<�����"�e�!������Q���XZ���cS���pܑo��0"��`�B��rf�a������PX�)ǡ�����������
�y��S������;<QE����ĥ
�9�풥>�i)2��$���w2�#k)��4�@�7'd�l!�Yl�������i"���b諘B���"M.֣�
7.)A��c8��c�k6�Z�XЖ��'&�_5�<U�$>.m�Y���}m�Y9�[4~���<���xѣ���f�F����H�+�V�y"�ǐ4,DZ�އ,S֮��ʁfhN�a�g<	�¦�I��ö~.�_瀀��2�k�M_#>G���>w o�� Bgd;��L!� X�X>3t!#i�뭁��<��L��ke���D�_$��S���"=��*Tf���/��]z�B�]-k"���v����q�)�OBf��'=<��3$�k[*=y���m]��Y*��L��XOAN�����j�lc����Т���U���9[�����XsY���Wa�5h��+4�<��g(đ�4&a!4}�$�ye�ud���>J[�����R�u�)t2�~��fm<������p?�����c��|b�:���w���F7%f£/^55�+�8�TeJdk*s�{�\F��~��݋��<G�S������1���0�����bڵc"V5R	A�����L��E�e��6wp3g�t��[7�·���>��98t���i��Z��OG�Y}ҫ�MQ�Q����]�4t�,e�C$.��&��'� �p���$�����_�*�"l�'z�{�M���>��{��ħ��O��+0Xu�X�m_��ȹ���)N�[����?�ŀ�#��[U�!�w��W˧x��7.O�BJ���l߿��1j��u.Y`Ux;��Q�>[���Ey�k���@��f�������Vիѧ;v��"q������y���N� �f�����Ee���Z��EE��J�Ws�3@U.9�������ҡ.�,th���s��r��<ЌR#��ɛ�O��;� ���(j]�b��IdJ�Z���J� n��-���fh����TB����KL�6{Cp�M��T�:�#K�7
0h�`B�ݝ��b��lL�}' �/1��㜢�=А>�l�����d���v�\.t��cB�7���3�H��M4�: ���W)��8��.0y�A��_�C�ż�s�w��b�ꝕ�!��p�r���	H����G�~$Օ�6�O�FYA�W ���εvK� �V�������v�7p4\��Q"���0�Qy�(F��������Ѕ��de�w�js��n�# UM5�'�8w˚ajj�U�T��]�E��7��.�zO}.�&��Hu�i�"N�&��.�+�3%2�`GYҏ�
G��ݠ`������ ���)�̯�������?x5o�rY�4��PaZ���'x��l�V���P��R��1������9�+}�$Im�����̙��ۋ�^t�QJT�O�D�����p�
S3�Q%!$��63��ݏ�����Ys�#��-1Y�ϛT.�i&����������reFo�^9��_y�R��,ݪ�5"��-���i��l�G�zcQ%�.'���(y�@��IR���:����D�,���QG#C%���u��ȾZ"ɉT�W;i��S�x���[y����O�]X�I����(~��U~�>-B]���I{~�^�c���c��ҁ?Q��l;��sD�>��_i!l���2��;�(�������N�|��m"�
��N�\2��8�:QPO4w��(���Q�}�9�N��Ak�P�����'��9|����Ѹ��m���?+�yP�I	)��<
n��y��������rɌ8����&��p&��jviCc��0T��*��д��ޥc,ૻ�n)>�Es�o5�X_K�f}ҥQm(��cj(�dc6_4��ֹ8�Cn���E��iR>�m��<��u�Y��7���j`Q�@B�ߎ[��UW;�P"�x�<t0��7rՄ�ȳ��<��0^(�b��$���]:{��H �<]n
)V>�
��z�%�S|�S���٬v����}�;��>��:[3~��N�N3�(�|{K^���t֌ ES�[�*G����t���c�]��hA��_Β��?�p&��Ҋ�^���%�5��*����5ݼDW�U��$�!aG�;�j��;��Q�ϭGZeԍ�|`!�D�O��Q�Iy��	�{Q8��M6�7Zn�rMi�or�X�n~:p�Ƹd���e��K��Z㾊��N�w�oa�@O>h����.�q�Ed�ZE�x L#��>0���3���e��7��h�?�P�nBtѩd��7Al��ЮH_�����0o���7E��U]��}�JOP�b�A,��9�O��F8�4ڗ���C����ɍZ�ُ��Q�8w��4��V�����ugMɗ6�$��g~���(���6��9K��_�/�xE�:0²q�"ɘq#�X�O�"q��v�� �1�6G�hC�-��4?[֗%X�ް(|=f@j�A��j>��L�m����W�+M�[�_aE��  �]��:����n���U�^j�|ȣ�Q�� ���c3�#���除�O����J��Dw��("��kM�Z�qL<�p>�L�f���ѣE@�Z^���`���h�����;w�|�w.c������W��AII��Vjǳ�3������O�L.-�F���av/\�N�[�c��nk6�ɟ{6h�����}���gֺ�!P,��p"�)ݺjQ��w���dϫ�x^h��EkD�٘q�K�Ş(���&���48��ز��w���>U^�(v���q-|t]�`�I�W"�NOjy�ҵ$��9Al�I��:��{~��*�S��?s�Ԍ�.ɐ���Z�E2��8��C�N��ӹ�)���<ru�$&��Z�0�k���'~�\î��,S��Tv���k!��&���l~�C�{���_\/~*]\"�8��taJ�����X<�̮��},z�Dq�mۣ)�1���B~���Gq�"���-���X���$u#a�U�V��fǎᒍS�s��B�u�`sk~�`�W%�XSD�?�=S:��sC���C�b#�n�L��2�'�{R8wnO	Ao�$�Q��+e�p�x|~|]�Pk)TS<�%=��Eh�Hږe�aؗ���=����=B���'[l�jUk�:�(Ԇe�(4�MF�}o8����������2�lvq��G�em�x�>��<���[�YȠQ��}3;�'�"Z�����1����=Y7О�3F�e0��X08e����"!�Ֆc��{U�'.�w��\�#�~�zL�ʐZ�e\�o��a�sG6E�4�4{Z��V*�����6: �����?�A*��Y�3�R��S^i8Lw>�h��t�����ݛ�����N�M<%+�q<�����n��� h�s���5F�WO�@�~�wϷ����M�g��A�سȸg6��꩷����0�?�a~%�X���������T��M�,�϶0��^�x��]gēJ��6�v7E¼h�̑�^�W�uF�A��W���!��{A,tnC3���[``��6�uq�O�Ƴf5~(��+V�O���'*��V@>;Bt�ʍZ�B<��>�~�s
JH��ź���ifL�|����I{G�a�	���n����ʒL��HkA(�b�˅V��:��$���3���g�8*�m2�,ub��Q�#�X���<��M�(p���Tp&p��:]�b); >�b�B���A$�Rl��m��}�C,W5_\a��ڲE�uLz���)�Yv?��2lj�Ht0a���੸-H����萢Ѭ������f,mi��>Q�]#۷�l}����Θ�LB��c��! sL����Q:(���Y$��RV�c�`Dh��V�eQC1)Ir^��+��̂c�\$�
�����N�֪r��-��D����3hJ��~cq�����t,k@#Qd�C}!Ǉd�L�֩��/��p�gŭ�;���8�D��?{�E�ym"�;�m��K��!��z^�o O�!�cH�W1x��L(罋xi�x�I���?Fo|h�O���H�h�FY�n��CPû�IO9U͇�� � ��'�7Q��O������"z�ć� '�(?�b1�w�j�=`=M�a;��na���2;������bv�H$��Å��=B�����<7���5�۱*2%3�'3�37��P�j�D󛵛<yE��Ӽ|&�g����d������<*��&�([�j����SҍAK��J��.��pI�q����/�硧;4�"���s�՝��Y�.��u���m^����m�7o@�Pﱄx����mC}���r��5���������>��.�*lV����pG��\c�����;��:�!�GgU�P>��`G%�0T��s54�����<���I������} ƶI�S����X"}��	���>s�l�5��io�VJ#^�ury
~�@X�y:���]Z�s`��큖{�&�`*�#z<�K~�!le�Z��j�?0$�1���Z��/����4�{���ia�$a\�
�����I�����N�:S,��A`�� �)��J�	d������q��^�c�F�<.?���J&>ZI|!�H�d��V���5�n�|̮���I݋�\%�W������#����������/��It���6���3��yVR݌:H����uL�y����l��<�s�A���=	X�["Q�u����z����IW���:.��j��3���D�'��o�Zw��`h�R[~앢����H&���#AF(��$�G��E��\�M�T=>���ۡ��׻)�]D2|?�wR���9dtis�j���~�#�M���7�]n��t�	��0�����W���Y!+�H[o�����O�A<���jn�ܡj\�&�kde��?��l{;1V�7�T%��N�ܣ�?Pe���J4k��J��c��*"���վؤHx�c7��/�t�'y gė]�Y�����~#���z�m \���r�\K��]_���6����$:�>��=�D�}�	amI�c���Q.����+�h�v�ol%�+Z�.���.0?�)wc�dMc%h�t��[�
�K[ H�T�b�u���fmKV-�Ți]��O2��BF|���صץq��1ӱ%��o�D�}��)�������R�Uu҆�uU���	gt�^�P�-��~\Z�I��¿�g�{s�ip��賆B�4��������Rw4��CcEWۡ�ʯ�z�a~��2��m8��@T�;r��]MkxG\���F�I��D��J�Ў�L�׸��{�����M֏�c\���-6��Gŷ�`��Kd�&/�km�*���:z�Yn�b	�r�\�~(��Qr�z����O����(���38��ӂ�A�^W�PSF��İڢ� �Hb6W���L,-�9�TU��L�P�5��/�|Y�ġ�T�货�7\k��>BK���y$u����8��j��qD���n̺u�Q������^�=��zV��?�zM�b���E��l���Ϻ�jZ�~�(��Sp���ě��������V����T�g��=���A�s�iM���k�aY���7�����
�7�6���N˞=��}jI�ܷ���^�k�zA�gcd�^Z�׈��"S��.�?_D���=~v�:��;���Z�H�|��&�'��г:�wN�0�I�DXGKb��u@; H���o�����kU�B�Q/��scB��ĕ��!���f���nJ�K*l!�:?j��Hy��};7lX�kh#�H/�p��q�z��Ro��&r��0��*�Y�X�dG��*WAPj�H�������z2�:�RTg|/����;"1kf��}΃)�k� 6�\�.p��������2��vL}iɔ�ݼ�	����{w��-��� ��p��@_�����g����_qk��ۛ+�'4κώKRJU��8�b��Y�8
l�!L�Ed��Uo�C�.���W��}��� Dѡ&��_\so��wȂE!71R�k
M����E��� cѨ���TW��B!-/�h0m3~���oU�5�TW�Z�n1�g�j	=��9��q�R�<J;<�d^_�M"a��1D�=�/<�;�����=�Td�̧卢xƨ8��^�w)�\}Q`���C��0I�V�I����O��߶yVo�t��o������H�����ݠ�Zˎ[=)���SIH�� Қ�قdY��-L�����L��!h�'��<��τ�k��QEg�>�/�CO�`X8��/'��!��E��'0�~�� �Lz�t[�-��,_Pe#Q�򺤃���� �]-E[�����.��/��=j�<�-D2��g=P��9]�A�g�ly���ڮkʎ�3�2p:���W��	d���גKT`[�m��s<���tZX����I����D�O�����VU��O�Y��=\4	�l�؍B"`Q�aY�Y+�J�X�)J1����X��������V�\�q��İ`�^����:<����AN�Od}���D����}d����5��X��p�j�1&\+�����P?��B�j
;Cw|�"fEJI���|8�Ͽ\������J����,P�B�v��S���q�aQ��"�������l���T�z����[�������L�f�ٯF��k���{�u��Q)=)z��q����TQD���@�}�B;�o��k��%�Y� z��ᇃC��r2�P*����t��$��Y�H�QW���Xr0�h�'�����m�W-{0�i���?�r �]�[#m���A��B$ViQ(l�q/�x���@޷(��;�Ȃ�a�s,�K~�)�-B=Ł����:�5���l����36��n
������kq�Pt����&j����V��%��*���r\}�&���@42��WL�V:��|�sރ�����?�2=~�G_Ga�ի0+`r�>���$�"��E��=`�<�6����S�DI�sV.U@ߏ�1����?E���Tn������"0z������#JE���cz�A���X=�}�2�$����������4��'�:�![���*ls=��"�Q����~�H ��H��>��ؿ�43�& �΢��ف#���;�.D����`)��B%��UQ7%so��������U>�Ȧ�ϑ�8�F�x�@�GGQp������F�1�h=@������������b�oc)�?���/�9�i"�-�w��eVB�p��+m
jҙ��>��\��B�#�F "l���!��6�;ٸQ{�c`> 3{
(�$���*�ς�h��aV�䱜���?���P�O\��ޙ�c�l������@���F���R���T�P�����3LR�|xA� f�P�Xq)�ƿ�"��//\���uK����H��>ߤ��>�7���322�����I\�{�N�"�n/q�|��a'H�1�=7�YĽ- ,�X6k��o�g�YM�n�wڟ[4�L�� $I=����?�όE��?�����q0oX�F?|��g�U�%�a�'�Y����$��"�{8����{��.C��d3@f�a�����p��K@��Df5��<:X���;�MƩ���1?ل*�3F^ON�?t�E�[�(!�p2Jdk�g11ñ�0�g�x�3�H�`���2쟦:s[z��)�IN�\��hXV�|ǃ��)�_Y�(��!�z�3�C���I@W�L�ӌ��~")D^Pgp��-ħB�a���̋*װ-.��e���2z#?�< �8|�],g3	��i1R37�H���f]�CS�9��W4/�	R��ےg��@(���QnZ�o���F׭�Ќ�E�&WeB�'J�yĬz���`��)�����L���m����r��=;]�P;��_	����{u�M����M�������ҭ��̓P J��t9��.	)�/0T"����ׂ����栎èΧ�酘�� ?�ś�in��k#½�M�ة����Z���^3�Jj��:�4k�U
�AETw>-�AE`u\!�]w:�}�u| ����[Đ���^����c�C�Q��:�z�Q��G�d�Eӡ�>���cO�Üe�gY��i�<ϔNE������Ɖ'�9�բ{�8��"]��3�b01+��~FE~g���YsF���;u���e�; ˽�b��|髰��)-�Rӡ^Ë50k�*QƆ�N�z��M�����L��<�tW\" ���/&y{�Z1�գ��ԋ�+V񘤾�I�k�Ĩ^UO��|���T*��A�m�jMz�]>�s�C�+�M[��r���n6�Z��[+�i�=�.���Ն�|]A�̹�@=d���?Ob){c���;ٌ�!C	�R�U�^�`���]�1�d��Z	{Y���}f:��`���h|��_�҄�[G%�!o��iP��>,n��a�r�H���#��&CkZ#���@��^�:��T�VvW*K���?Ri��$g� zw�\[��4RR:��!�K.?����3�;����}��X����g��8��#�3&m_Z�w)�h�#��ϭ��C2	��w�
N���������a�v^D�kz@�k����b�$�5���/PdUD��x����N8���!S�ӟ~1l�Fy����з��S	Q���d�m�����ͫ/l^IF�&h�0�d�[�
�<����TƔ�hq�V� qQ��b:Sf)�&Q��T��m�xb�!��~dM&2]�ϓ��s�	�g�L�A׎=ҿ]��ߔ��ō��YaM��迳�N��w�%.�yVr��i�jI;f�+��JQ(_n�e�}����NF.w��a,#�sEvF��?1���0}�P(�NWpV�L��������/2Kj�ƹ"�j�W*��n�K�C�N�J�}r��p���8�AFʯ�R�GƵ�"�oKkv� p�}�� bַ�1^>�H�����mirEO�8�0>�����0ۨ��PV`C8J����>�����h�o��o%��FR��@�(<���֞L�\���(kN��f��q��_����E��;�s	@Hvoo�U~�U���5��G��p*k{ger����q�۵�����K��<��Fu�D�!z�Y����̪�;B��k�{=�w��-�����bơ�����R����s�t#o]Bؒ8�ȬXv�#z�-�(���zG�+�j��b�F���-��m�v��(M%�mf�H������o�AD��?f�F��?����7^C��:��8
x�bשB�ج��O�s��5~M��Ȇ�kO�zԒ�Rk��m�?���x>�j���1)����&N<=��!C �5���:��ӫ@�NS�(;0ȁ�62�b�w��7��L[!`�ю9Pk����3N;��ʈ3`�	*�d�J{781$>�`�v��h)��?�{�S�rv�̿�@�����7�
�Q��.����(a�Z�tmf�3���[�/�F�V��^IP�i�uT4U?��,�r����M����$��ύ�J�)!�ƌ�?q��s�0I/b�/ΞLp��'|��y(�F�P�X�~�T\�������F�4���4�F!��n��d�+���a�>M��XK���ǁPCkl�u�g�!�Fu�H>z/���L����Ђ��ۅ�,�C�M<�ʮ�+�z���K	DJ�x\����e^�92�tDGŬ��a-�<U���2�.�t}�Tn�T(ŗLԯ�G�Gw�i�4�J*�����6%�%P0B-�tS� �t���58$AO3�d�'.O+cz�3�1����v\�����C?ua˲�+7U��)��A������H��?��BL]����n�;�����x}W,��4R�e/݀B�	����3Ed���˞:"J&t���ь_Q���n��!&��y��2&<�������#:�R�k�Q���(�4��i��ɥ6��h��2���a��C���7f3u�؞~�2�3@�|�e�X�Q��^a6Y6�E�����^���+�Q3�1T�����#)j\�JV���̃��u�iZ�������5�A��6��4����~Jp��9g�ޖ�9�_%+ŭG�|@�e݁b?��{>�7��G!6�H��\I��?��q):�L�S����4��-'��O����,��3͌Z;\���`�OA�z��|.��<���g�/��r�)`˨2���&�m�j��>] @\֡���gO�/��{>�k�_���-�#z	���ǯFГ١���m�����b����
J�L�oH�	����S�0��OO���%��y�^��ӎ��C��T����ė�ܔ'�L��S�D~��V9	3;ŜF�
���� g�J7g���)}����|E�!�|����1�� C��@��J۰O�\��]��߻��|Lϭ����ӕVr$���{
!ZLyS%�4���Y]�˱��d�p'�6k�~��4�Yx�9�k�d�Q�0���	J�(���7H�,@��R�t�����F�4�5}�&㙿�?�{��RZ�G�wK��Ԙ���:����[��9����q��mr;pB���9nl�� �l?���3��)V�?�<�U`%{1	���8~:#����6��\������c�E^��~��\}2
��J^��zz�B�PQ���2��Z�B��cS�~��#f��u��C��s��v;�,Ϧ�,&j>�E#b6�%�K	�u_ۘ��8���������tc��(SOo����������\��1w����7z+��j\YD7D�5a�F�+�Ѕ��eLܥ0�BT�*�������\���+Ȗa�D`��x,����iz��dd_�t��N/���(�2�Tƾ[ �!'q�S�%��<+�319�R4��z�k*�'I(�*�81�ݿY&����cK0���#�dw�j�wm;�Q5.��(��dG�e{3���<�n���Q/@El\h)�,��|o�����c]�Ί���Yx1s3��F߱l��+Rϼ��l5���P�՗���O2�5�a�;Hb���V�)�,9`���9Jڛ�
=UZ.��9;w��/sݻeg��J'�Ls��h��*}����r=:��*EX� 
��l�=k!l�>~s%��e%/O6��[�@}�)�=�v�nQ
�(�l��Ǔ-���.�+z�v�?�QA/kXW7��.�M�D�e�:��p�P3T�{���cG�rE�</d�H�X��b�1
�i���knC�~��d�5j"��|���{ц�Z�p8>��aH�)z�=a_}�_��nm�e1�4���%@[Ry�V���V>?.��K�T�S�T��~E�Z���V��D�
�|Vq
��z�a
���!q�k޽)������{e�Pn\�m�=����bdn�>p�Ag���K�X������u��d��[Z<�T���������$��u��h�?5�Z�N:�R��Ⱦ��^� � ��pZhe�������Y�q}�b�)y��Pw���hŻ��7AO��iJ����u���
�s5��9ٳN+|C��J���
���8�C��]VYx����Oh�`1>�"�O�����/g�1�B������UWE��N�4�����x BR�8��I|J;#ec���i<8X����!�;� f�m[�g��{vG�p����rQ�#�!-��"i����|{��O>f:�|�w<�ń� ���T&�hC
Tb�nO�U{�wXL>��G}���6�]F������F�B6�AoV0�q4X�wb�3j';���#�����zxf�x�+i�G���	�PXtNꥇ͉rJŃI�w��|���{�s�\�y-Z�i��c߹'
GP�� �q~�>���QOJ�Q�NI6�_��z�ge
��,����'4�(��G�+��[�}G�;�r%�%O9�E#�
�|�C�^��4Ӧ����������G�B�,��4h�	�l?��RoG�����{6r[<H/D:|ֺ�'��wN���%�hci�ճ�G��_�Z���(Q��`��s�K���E^������3)dI��,!������ѭ��5D�e6���Y-��v���{kƱ8ju|z��y+��9�(��b��%��ؔ]�+!v���I��tT���@��Ϣ�!�c�^I}���s�a�]/�:�=���n���}�[
���h���+������\�����������I6��V��^EZ��_^��C�;��a8�~�V\����f{�f*~��<nj�g�D�H5>_ �*q�|��}�'��\-5`�K�m�/'-�m��|^/�H��{*�Ep�����b�/�v+x4D"���k�7~��Z���d�5ՏJ[O��B'�8�O9��������h?����V'�O��qN3\��+L���i0�@����<�X$�H�F}�^�����=�#J�`V�;m`y0�T���ю�?�'4$�Ӭ�I0�$A�����&���%���t;.��ޮ��I/n�*]��>��c�`�[e����
���z����/�DA��ٙV�t���}���`^|�O�%z;H*ry.�H�g�q:�s�!��h%\Ɵ���z�Y)��m�y��&����Ԃ�!�nn�/@��d��� �X�Os�a��-����S�����_S��f��hSA��3���B\]zh�*b:�z\r2�o%�+tfΨ�$xM�祄�^ҤI@�����,~��ކv����)�.o'�h�� OAD�H����d7f�Q:=u�����٭�N�[~����:��|O�?�Y�����eDhJ�T��"|)y��}S�m�����^s����;h?X�3]BLX��C�Y���-�9���v	��3Y��N��ᝐ3����t�mH��~��E�1��y6��i�4d۵�Ϋ�$k�G}xq1J�Hu��B	��3ZKl�������0��lj�.��H�5���:�F{��j�^ �@�ZHAҟG�������;m���٪���{�,�.�vg�%��*���e���4�������)��;�{���s����[���x!N����k�k��.8�:��(l�PB���̙;Ȕ�c`F;�UgԠt�M+�m�ִ��2��]��Z�Eq�3I�QJb�+�Io˞�z����N��;Ю���ڦ�2�~�b��GP�;ה3����QE�B����80�dΚ*��.��M�u}M�I�<9�c3	�~6�9w���g?�ӎf��瑃�G�fd�=�:�.���2���i%�ccA�#YTT��]	%���7�0�N��TyCW5R	d��_��t���_�P9;��T�ˇ���75"����;�S`�r�o?��X�����p}�3v���=���53�=M/��U�Ξ��fb�����M�W����piBx���۲�X�a����{���l(%�
�d�|˶cPȝo���!�E?m#������0�8��S^Ƨ6�o�̺�y�U��)P��*5��^3&J�?�����Y�y���1��χ��lj��� ������O�.���t����;Hg�G�Q~|�R~f6�_����:_ZTF�Cĵ���
�#�ȯ�0����'"׶Q[�Y8jw37��ɹ#��]������D��'Κ�TQ5)�P?9J�\E�.3`^nt����[Ru�_p�~��I!V[��{{Cc�ζ'��ݕ�����C��$^�(��2!"���3K��#�Rv�25v$��H�,��`B����C�_�z��C��̦��M�e�B���A�ǃVIa	��
>��)/�p8���T����p�'ˍ&	��Կ�(��Y#�[5�E�.��UJ	�F�:����Ty���e[�78��2�'+j���'��߁Xy^�+_♑̪�0�K#a�[�&q�
Y��i&niroK3��
�[���^'����EP�p�B祿9σ�pS�>~G.@�Hul���Q��/��(�?���u4A��}Z���H���>��1|��=}*��l�4f{��W��'�/�m���_Nu܏�{a�Um�����S~�g~��T0���_0��sJ�Mdg �[�_�K�zF'����]�o��+K�҇x;�b� �f}�$��מ�ӎ���^��s;4��ߓpL�� RvZ9�M�V��5����,��w�F�W�58|�
�d;�#���6Xdho��ԎŌmH�j��\��@���)*[���e���x4Um���8��_�d��h�鑈q��\K8����-u���퓢�-Ph�-������M|֮�PNo&Ke��i\qT�!�E�o���͗���N���=�
Tz��0� C P��;|�$��3J�?`�$^U反Զ�dJ{�V��I��M�A�n��{n�ڽp��IP`��S�ES���p�؟ϒ�+p�˘�l��u>�獆��_���U�n���vZ]U���b��H���
H����V�!Yo}Rz�޼Y�AI��V�֙���8eA$Kk���R�gmaxL�'&E�9�S�u��XI�1� tJN\9��@]n��V����ؘ} q�kl�`��� ̶5�K>fn���wkl�����+&s��],��"��]���1��Vۖ)`��bUo;;���W���Jk*�z�G��%HLS�@D� ��Cy����1'�E��˲�����qo�r-�� �^u���7®�]�J^'�.~ٸ�ӳ[�(s�.�� u"v7�ٍy���P�g� K�5�Ь��_�O0yt�pQMr�?����镐���R�3�cfO�]����|����e�%NЙ�o���7^ٺ10Q��Pn����tT�5\��I`h�\
���@\{���PB�|����_�3+����N���*�k^3D���!s
�\�c����ȴ�f�]�+Qퟆ0G\�D�4�N�P*K`eI�q��s�#�
�A��R��߽PW��s���E�4�o)��	�c#��Ԙ<��2)�e<���;p��
��mʮzM��U9�"�K�Q-�u
;'|��&�x���Eϲ$\ѿ ��/=�,���}qN��u<���_��b̼�wp�?c�!te�7t�&��'+��i"�k��@]-��r�SoC�#\fٵ@�b��F�7{�tKU���S�j�ۃ���b��z��Y�w�t߂G,�T�G�<�m��D��&����x��i�̿�:��fIteIn֓�������$�J.���5U+O��%���E���X��<\鷨�����ҕ4�R���7�o��	�[\��eλ���>\#��ܹ�� M�gz�W�[��+��!	:���I�v�������
�'v�����-�⪓���3Q�:âޙ�i�6$�"倥r�pZ����Y�.�v�l2D�����|U?�L�Ot�_D�X5�dk�'�^�dBa�S^�x����>}׮��r�s��*^�$|�z�y:�8b�*��v����9CY�4%K,s�>v���&Դ�O�<�T���;ng��Znx�6���8�j�6�<e�Ղ?��!�����9�.��u�_���y�ձS`F�D�aM~����(]�I�������8����~��c�1Ŷ�0tB^=2�Ge��Sw���d�BgP=3�%�lk(Φ�FЂ�[�^�����f�%S�K?�����>���W.���]�	�쁲�9��[��s����v���q?�c�S؊#|W���NFH7n�Q)[غk���I.-eO�%H@�1Q��WB���M���u
h���	~?U�x��݇���@�����2г�!�H�r}Qq|�RC?���Rs�c��8�� (uj�}Y�)t\�r{-)=F72獞Y�do�y7����#��|�����b��K�_�kz`�52�E"�'Zq�=*H�Yِ6��$��l�k̗=œA�K��A���N��4��Ƌ�j�0ro��}�����1ˎ�7�~ٻ�.�eȋ�_���~ ��C��3r�B����Bl�\��� R��]�n�T��Z�@.�۶��X�s�+ɥq/��'�h��$׺�����`�ޠ.��J���R������ʦ!g�9EqI�K��o\i^p�vs4�]#Pw� �����X`׍�?JM��)�A)%t{���W��)2]��q��ܭ%���x{7��a-���\��#F^!6m�]��Be_��+�<n�� ؝ȘH�D�T�W��K��r ��0.Q�oxh�e�\}�':Ы���=Y�2��������A�h�]x�/����c;/�i�1;����2S[�Y�`��J��&��2�P<�̸�H�h�(���iD_OP�ͱ8��ea��"9� ����,c�j�<�|��<�=·wA�`(c0��ڔ�G�.��ݬ�W U�O���d!O?���}7���K�^V߭>1$T���D���|l$������N�{�Uh?�c�f����[9p�҅_������� ��,2�r�)���Oz�T����Sp1�󑏵r�~���S%x�t�j>��/��v`�)� �Ԯ�?�J�h��U1�m4j?���$;��/\|������o
f�"���}ֶ7��p�k��zY�P;B��:�,�el�6��X|�,f�����G�7s�DK�H�˖1҅��1��Npz��G����E-�O9+B��A$��t�i��k҆<aU'G����{�FH��	���tA����M�[g=�N��8�q�c��-Iy�GF�����ZQ��rzܓt�x������F2	 ̋)i�����VA�����2w?�Db��d����dR�
�������â;p��L�x��T����_�VWY:"� QP����*�-u%�Ԝ>��Āno�-���OF�Rs�z����'���ؙY*��lν��/T��������8yf��0 ��F�_�Y�t�7Ul�F��{/C�̀oX�F5�hs�
�B�H��L���MYp��]���o%#��s������cϬ�+R.�͡S}�K~�|���1���S���˄Ф�����McF_k��V��i^61nb��=pE<�j3�䕱�$�6�}X��c��`�6�]�3Orx_�Y[f�j����{L�?%%�/Ut��[m��W~;�	���J�s�"�ʆY}�5��{�����⁧��P4����ckUWs�|,��D/PkU�A������F���
��ll�ͻ|�,��Ω�E{��OM��`"cd��#>�"	���9@!��_�?�ԟt��ĭM|�=rV6F�	WP��]2�[*��t��FO�&�d-�%���W;�`�A�ň����l�d<��֨䁜�{;/~��׳"{3�r�6����E#3�-�C/��y�� �߃цe�:�l]0���A2��*�����Թ����yXM��,��(���탺P�h�`y�͇nA#n\>�2I@���~�br[	dcm��V<�y���F�1rD��;=�e�`���ҞZ�|��dO�*TV�>��#dR}�������j�P��M7t�bw�Y]��q��ڪyf��,��i&�.L��Uְn[%C^Vx*�H�ԑ�LS���zJ�Z�\#��L��(��28G�~vc6�
R��ŉc!�R���Þ�������a�+i�ɤ�v�{aZY�һ�P�s=2hg<��	�2
���uJu*����`�Ѭ�hK���ѻ�;h}�	�e�D�U]K�/':!�G�.�!� {�����D2�]���Sˑ���a�wsS��|%l��RQ��rx�+��W�-�b酫M�|K�	����5��MRQjB!Ioz���}��)pa���n�Èa�wS��F�GH������-]��d�VP�@�i�����HE���G9`��
 ݁!������j��F@G�w��lz���d15Fv��{�S  I�����J�խ l����l��hE�S���������Dn_�Z���}��t
nF�N�!Χ{'�"M��f�j=���0��WJ�����N�T�9����8o��̈��މ�w�K���5�����ڰ��G�ak)ˉ`��f���F�V6u�'n�*�g�2U�D|� ��0CS����nϯ�]f\��S(�H/��X�iǈINC��^/��c��/�n8޿3��M)��t��t�Vܶ~x?�z��u������9b)��i+���FmW�G�6Rv�x/fD�m/a���h<�nH��c8?���gK��� ��e"�\b�oh���t$�W��_5�Z�?��ze��A�
��ړ�=c%��z��i��L<W�#ᩤ u%8ȗ>�Y4ZG�2��c��0G�ig
�m�;�m���-֜an�ԇ�?�[��
��up������F��J���Ἀc�Fj����X��$�,
}-(P-6���Wr^l�2�A5�X��<�Gw~�Q�|�RU�p[�����GR���'���[��q4��?U��wA�M�]�؉̄?��);�n� h�G���k�q�H哌1�K2ؓ�'6~�t1�K<��cw�ҎN�'|�
�{;����k�JM/��]��L�[���ٮNc�"FRS�4��q�RXY�-(����]�3���i+>qԜdT�|O�B��c���WX�o�73�:z��qSej�f��Kׯ����OF�1����F�МgIo�����SC��^��U���K�e��se�"0h��g�d���<��2��N*��\�g�)PD�^�?*b}2]P����v�[py7\/�k�@����<8��y�a�! �f%Y4�0�4L@�A����vv=mA���u�MK��-��s�V
�;l��ͯT�~Da����b�$ʃ�J�4���4geԕE������+s��<�٢V�K�hrL��	�w���W�cy�ɴ�b	l�#:B��?|����-�;�T(\�w�%�T�E1�K�
�z��[U���7�Ν`�.KZ��+%��(�,a�QMd��:B!Kjd�5rI��n

ő*L��b�+l�	E憙�8L)���2�9��]��*�*tGAJ�uG&�pVA���YN3R�/r��w?[�����s2��ao�(��-�K�`ﻄ�b�a�9,O#���-E)9�U�OI�
�4�7�C:ա%���m&|����&Ѽ��"��*�?T�'��^S$���+p�N�h���CGk�ъ�)���?�Z�#q���C��7dLI�~$m�0f�I!H�\r����D�X�D�����P�9��������?8�C�vV�7>�ط)ܶ=���&w����+֡��EC�`����q�]k�$t�u��N���u�~���L��&8vtr�C�I)�"Lh�k��a4������g|T]ս�
S����Ear��&���b �J:,���N�"S�H�RE�qY*�W��|u�gr�%yXohf�}���&��4�N.f��/���C�����.�L}�؊�������䧰��&��y��}������<���Զ�y�����������D�n��GC)Ǆ聹\��L4J��{[n+;���M�v[����v���g܏
�%���	� !g�z��������̞����̱1�g��e�S��ϹDY�9by�{x���#�EF%4�D������DP�ծ����ޛH�*q]����C��v�H���+5�_�1+�N5v���� �@6�=��1�o���W	v]z��i�"�#V�}��\F��YӁ{�#��zfڍ
�-�ʧ�JRF�p�tv��hO��ӊ���8�����d_Mc�}D�Ӌ�� 2Aq��5I"U����C~$oj��
)t��g�2Q�T�Ć��CU���
���n�2�f|�tљȾ��cӚ��ogpA�j�-rkRu� ���>X���`�%���(��ުV����=�R.��,���P�{�f�u����I��0��m1��� R���0�H�o(���.�Փݿ��=�7�.�Q_��{��ER� �`4�RW�R��I�1Yu�nZ��|X�D7�d�,eBR��Ԥ�s���H��a)/��
��k���&$n���J'"Ԭ�wCXB�'���6��H�R��bG��|Me�ғ��Ǹ����>"��p��b�.,�t��g����;��I	$�-k��k�n0875I� ͡�$)ɂ�x���X�����P'M*���M8����1b��X;j���yZ���@�0����N�$�ED�b�"]R���	�����K�W�M��n����pm̼Cj���4��R��jI@-��"�R��^�x����m��$�؀�[l �}�����@c$�_i��[�
rHM�9iƏf^_�'����8��Z��
��^߯�X��%���y;1�oTՉ8�V3{��Mg�����hOF�x���~ܖRu�eg�"���v}�q05p�JW��n���9+�������C����>>���[�����Ɂ�}�U%��`�
r�@fN I��i��c2�Ia-]�.l����R�����?�fL������0��q�q���O��TM�AL��7G�]�^ڀ��
����PkIw�S�F����=s�2�&Nn��!�Z�Wқ���c�l�?\�a0�(��✉�oq��6�	�`P��<�&aqLܮ�=�,+�T�C�5 ���K8'���!)4#e�flg�ie���|A�Ǥ�Aɷ��o���:�nۮ�{���� �L�P��%�ʌ��>TK�k� �Q��0�D���5S�_Zt;.�6J�d#���;̲9w��3�)|$�d�4�dٍ�^�Ad�: �x96�&�4X�@�a�r�[��s��'^�Nڙ�$pũ�M�x{��_8�����F��Fx�͜���ooat�۸��A�ȸ����L�Ĕ����97�}��&�-�G�q�~z09ًٖ��	����%֗5t���kpH7���w���1�[	~d��k�Ip6߯F\n"��,��	��2��z7dR���C�u�R���{���NmX7������B�T(���3&v�d���TT��I���Cy����Ǌ�&sO�p��)����6�I����Ⱦ ����(mO3�c��3�ĥ>=�] I��(���Q��;��y�&�
fBt��)2�o�Lv���ڽpN���ӥbW�����-r�	�ۓ��-�Pv<Ѣ�<R�X?*8�_8��zz@�]���^*���)�&n��BdE/�@\��s_l��s�嘁5�Qm���_����zIRC��u�b�]:�f�뗷_�'�a+�ʺ�W
������1� O�S/�E�j)v����n��S�HI[#\1�z�6N��N�R�>�u��IK�
�����&�io��6q���V���D4����j�]�W�Im^�a6��#��d��R��h	/Q�vУ�]�e4/_�˿pws9L��۴���x�&Wh�N����ʣi�`8��F5.G<���f�Z >�{u����t*/_����ꅼ�:d$?X����(�&�<���3�����J��dն�1�jz#�Tif:�ٕe(����� v�������[Hoݦ�	Nv�o���$��ן�p�p3aP���e|���XK��6Ԧ�5�����\+���Z������P�zա�P���~P��� A,m������(�^vG��H�N�7�pG�=�ӗ� �d�5���J�#���V��<v�3�|����4����ĕR<g$��
ȫ]��݃��ʟ���]n�O�ް���x�)����`<TƘ�&���X�=�&���<
"����ʌs�M���UT�w�� ��R{�kA�s�Z���'���� ���R#_� !��Ҥ2Q�H�B+b���@����ʑ�X���@�t4W����A��if����X���tn�����])Ba(��4�w�Ol��gZ�J>��/S*�����6�2�M�-Nrx���M-��4�e"H���U��3��)ޤ���=�o�08��E�}ڱl]y8B�������ذ����@�<���ƻ�(F!�$�����R$�j/y�R��hM: �Vd�+� �d?#4��n<���X�ak��#�3-��w(<�\Di��sQ��u?Xהm���h��?:�U���b=c��ӡ�y:X�����r�	!��t�bLT� ϙ��o��Q5����~}�8!v
վ�N���)�Ļ�΀ciʎ��0=ĸZ|Y�%��ԛF����̎���%ߢ�zIU�oЦ�K��W����!/���e�]�zW�I�U�?�ˏ1��,E���5�d1��C���(�B@7m�e�s�W)m8�/ʖ�@�?�
��O�qAZ"In�y�����G�7e'4��zbw��"�y�x��8��X|g s�/�N�;��A��yP�i~V>C+���X@�����4���� �7>W���F,_���95V��?]z��Xr��E�E���v!�&�w��ӹ�g�LF��F߇�}08��Y��)���������Pz������|c�I:n�� U�S�,��}�c{��2A�PU͋����aQK�$��^Ċ�Z҇�����e��<�����ڇ\��Ɯ��v���F�#�0p�̤&~��(C�|��x	��R�j��Zc|�%|�u���-B�8i��Q�#���8��*C=�D	%�f2�r�j�x�C��Yao.���W[:�L�qd(������ě���鼢��~��^�X���h�v)
��
�;����mF���a*��:Ha�8r4�3B�/X_�
jF�2��Yî1]��F�Ū��Y@�ᤢ}�5e�ɛ��j�AT)��lI`�u��u3ch����+z�%?�/�6U��CEB��e������Y�ʗ�1�JC
L�7���.&��8��"�c�����9E$ϠJ�Iф�0�@��i�n�xZJ����Э�1���X*y���h
�N.4t;M��ru���h�V��
f
+�ʌoy:�w������fj���=oΏ�|9*P����ϟJ|W]6��{��Ր����c��|Q��z;���g�_����De���$��h�v��+U�w\�e6�ʤ8Ŝ0X9�jR�PiVo��Օ�'�E�6͋O��/��{E���س�B 1㜎j��=h�TZ��uFsz�ufs?�o��N*§%	�h��ԟ�x/�$��CX�X
��+�ѫ)�4��)�,QJ��.��9� G������ȋP�G��V���c߶ TM�r�mwg$�*�I��?�P�V��^}~���>�v�|J��G�
=��,2�H�j�|%2G�?f<�� .�F$�k�I���c6�Y��5���P�ٻ��>����h�[+��Њ�?�*H8���8��9p_U[��j�IW����ctz��V�AW�<��t%��H��!��4��#��q�x�4�و��ü>}{�>���7˳e�>��G��T����6�!3ш���#>?E�E0ǎ��@�f}�9��t������]^2�T�e�����V) �2N8�/���~��?�l �#DC�����2��GC����b~>�}�M�؏~��$Lϓ�h4L7����E�8C0,��@�w������Xc�4�p<p��-���2V�[�<��ߤ�P�j� ���zf�U�e���ѕ������ku��
�v����&���{Q"���v�YJ��w��G��!*�S%�7���R�����I�L�����T=V�o[��,=�^�L�_ĺ�lP�S�ҷ�C��F����3�ާ�V��E��̂�Ӕg-�&�Ndt��,k����S���T�������2p �Z�d�s]3tx���5w`@'��W
��Qgv3`\-���2狎�B�[�C�����R1���+�2 D^~��?14p�џ�@�wC�Y��$W�3ucmt�i?�,��T�|d�0*{Ax�`���P�=i;�ȵC��L50��9��j�2�ν��j	;���FY�$��J�A�~k7�唞�0��Th�_Z����;��t-�	T��Hk���Dw���o(��i<�́uPFq�cO��&Z3(-},o���A���ȹ�$l|�Z�`Ȳf)�C9`.�9O���W��K�|c@�|h $�������%�[�mq�V��'Z���Х�B�-b�_]�c�S��:��o�H~�I�fÊǢgϏ��9��A-�U�� �u�UD3HY�d�_��\n��X�����
��K4�ǁا���]N�r�}u��ޘ'RKm�G��:tb�`�����x���׿�7?Y8+m���\ؼ~���ԛ�$9@$y�+���;Q��Ѣ7�K�}ϸޡ�-��ݞ�p	n"�S�)W�R�^S�Ό���5��d	����w*���4A:Us�#��@���}�Nͭ.0\����fԣ�xT���Q8���{�-}I�4_F�6�晼��D�Y��9N�i��ztY��V��?����2�ٻ��zŐB6}Giŕ��x%D�1���&��l������0���HN�2��3"����e��%����6K��(f�6�!��K�9߆J��S)���`5�g����k��p�����G��u�6\��i-�:�+��V�A����?��\,5��	�L���h��Ͻ=7V��1��^��@��So�2���+��7�~F�=�4R��h�����O�g�W�;�К+�s	L$�[��l>]���v��7�kl5PD��d�ۻ��9o�����E�L�}��M3i;�ӳ��[��(��o"�D�Y�w��:����٦ۅ�'���2#7A�ߧ,nH��?����(p��Hh�B?��T��w'���*�&��C�jE.cպ��u�CN�Gp��!U?��~���((��v���Yunj��v^1t�d}�HA+*�Qf8@�񝑊��sZ ��#�y[��M<����L� ԉ�U�*�r��_��j�G֑2�P%��\
]Y��á@��ǂ���o�W��'��?)��������D��'X�k���œ�hC�su��%/��o�T���}4%n���7��li8�T=_�Ě+t5�0����&�9_�z����_4����)���r�4D ����X���./�x�W�����6�P=g^4Z���D�K���)Ц��z
J���i�w+�]��&�#Uy�٠jJu�k�D}�ύQ�ma>qo�"ì��,�ovg
u�?
��ɫ}K���Q��'|�a�<U�t��r욢�h��W5�p�>*��R7��gm�U�o���{�,0ƅE�>���􏂚�"���M�r{�	���H�>3��2�3?�F�?��>W�%�J������î���:��nو�M���6�w`w�8����F86a�kE�H��E���6��Nq?E4�7�7�P��j��΀��ݚw@ht�3��x�x��>	���L*��9����`�����[��-��觅�N	�P,�Ӑ$`�g�9�$_�R��Fc��$�U\X	�����\����y�jc��w�[�
R�" @T��������$�&� S��s�KH_��c �d�oVkg�Q��&�pN0H���^�Vi��:��N��U)�w����k�� c��3�����<��fG���Y��xH�|�g�z�7$ �5��_VU�0�Yd�gp��K� @>�=y&�#�]�jjD��ø�ٞ������bF�։�w!�����0-�f���t�S"�Oߌ�]e4`Ź��`��}U)s�^Y���m�n"N��@��_���A����7As\���������'�g��֒��w�S]5
M�������ֵ%����_
����dS���k�"�>������E��������8����/�ʃ��GԻ�ҘnDi��q�e4 u+�˓�i]�s�j%����]~�����`��&l�~�ö����𠩮3AG�A(^�S�H��Z���1�i,�C�x9[M�7���0�W����&��^���P����S+Z?�?U�=��L=4亮�����"���gz&���_c���hov�Å]�2�Y�[�\���&��V|���Մ��P���B��*s.lB&Cӛչ�ۗ���/�r��޿}2g�u<�-ȭg�HS#�JM��K�}��Mړ9�/�����*�7':�잟',��^!��tL�|$բ���s(	������z���>z�F�%�;�+�!�pn)K5x1�G5D�C�kZA�	9��NTn��`E����=ɟ'bHc.@��ϗ$}?t��k+���@<�^C"�1pg�iV0O�|*���u^���m?վ��u�HR�@rW��}��Ɣ�hOj�u�"���O���-<Ͱ���6��\�$�Wr�t�g��A���+�'���u��+�44�L��8�'��(��:+�k��'�қ��)D)\�Pp�Z���K6Z/)�'�����ֳ�s�q������wɭXu���^�h&.=c��Fځ��k\�=Q�ԩ�w�Q�?�:,_�"�L�N�"�Z���#�OWN�Js�K�DG���,]����^���앫�o�c�<��m��P&�F�$�,(��1�~��W8I�"mM��X𭱬?����2�"�������ӝ�#_��L��o4>ޟ�C��-v75�q�n	0����$��p�'�X�v��������J���ȝ��d5�4\�Q�[�ܥM/$��O��[�t�[P`YyH�O� V�������d���ib����fJ�BԦ.%F^�P
��)��#6�M����+�4"Bܸ�+>���!vu]?�k]��B��(����7�qR�Z�i"H�ؤ��tz�8����W�U�8�-߁4�֩��$ ��+ۢM4sL�?�#��Nr�����_�%���M����`�6���*��S��ʃ0�a���_�5Ho�s:e����~;v�^�=����҇����5�i�����?&��?="�")�n(O�}z�!n��N��T�`�9�f��)�fׇ�IW>׽�14�Ă�7�qL�?"rA�8�:j��^��r�E�Iΰ�]�{e~��������N<¯�N2K���a6�!x�u�)�����o��=��g��a�?���Z�/����8�
6��,�b!ZضU���d���t��RR��y\o�X.�YDEY��������ҨX��:����2�3�0c+��ZHE[;W�8��hc g����NB2���W�V�����M}C�\��Ƽ�@;<^٦��c8zS�vl�����FC��h�k�6|���/3�8Hcp�@�����'�v=&z.:ND�0�� �/�(A)\���t+��nw�RKbɭ���@v��h�p��|A
Ƣ0�̓��D��� #񌰶{�X���y��/��P����+���Q����������iZѧ����I� K{|���E���^!/����f!a�}ջ�BU�����t�i�UG�8�4f��7��d!�Y"� �h�&���3N�	Na0�a�߆�>6�$�=e"�3n��g�{����>���--����5�n�ٴ���p�N��Ĉg��;K@|��C�z*��a��x/�	|���0̛Ϻ�\�)O�fe���\ �#�7I1��W�sS��"�Aj(�����q>�vK��r�1�Z���co^o��\&�{Ɔ��C��&'�&��Y$Z��sCz&�U���?��&�3��@#�&i���۷m�w�Vˬ�@=�jj�5�������r��Vk02D�b���<�f��cK��#U��/���:��=a?�̩���ݱۓՑh|:��O-��؏$Z�Or�z���R�����N�x�&�m3�4ݳ��!G�hI�d&�!�$n�h�<����K�d�n�G<H�Ch��h�T /v���L�l|{��qNh���D������0'K5��#	jlLȿ崙�R� +��K���.��mJ9��E,^�MJ?���~�ׅ���r�&� �+��W)��)�*u H	6�܍���c`ѿ)�ۊO�˅�j]�]i�5��~�ra�g�3πD�x� �����$��b_,uW�=(�'z�Q��3$��ќ�%)5�����21�"�'t��}ý��!�1^�1Ps>�X�K���^ ��ڜ�ce�hUA����N,��h�H��S�7��Z*b	2�۵��\I|��`�\ye�[�1����@��h���-�"�/��%���E�ru�Z�{�x>��B��C�%tԌ^����x���r��P �o��5�����?N8���lȨ�����iA!!�hE�G`X�ιI{�Ch?'$18�?�yƼH!�}P�lw�D�.Z���+��*�?n*Zۗt3-��S���z2��
1��T���	'S<�'���@�N�R|
0[˚��d�=�����2#� C�1�����
F��[�MQ�`Fʦ�!��ɪ`�4����Js~��0����@��>����0����2�!\M�ؐ�3X~�.%��
�
ϡ���"Lfd>�Ԅl\�J�cʙ̠��zm=�l(>}Ҍ���C.��ϥ�������o@ <i����}�8C~��C��bg����3	Х�c�������Ib!8����85�+R%"�CJP���=��	�@zJ�ߐ�; ���J	��Ʃ���]���>c����ds$�:��Ŷ�[Al���ݗ�V^�裂�+����D�M�禶)��*P�Q�E͡�[^ �R�B;uK풎E�����X�h�t���;)���1��\�$�� ��ͶN;��'O��v!�")#�=�E�}�x;)�e�U��B�”�R�nHmx�X��iW�1]`�vMB����{zIߠ9���3�շ�+�gz�a�ޫoU�ݠa訅�Z�Db�:R��-󼜓)�l��-g��:��G�B ���s�@5�%P�������4��]�`b���B���`R}*������S�����pH�խ��$�q\�3����e�O�T��| �o��%z���of��BC��	*����g;J�Y��3[���w�ל[�S��۶�)v�Ԁ��뎙!zI�`��3���na��QL�KdzP�!O�9��"���s�5c	������^�'��J��q�>	D�~�	1E��_:�D(Twa���u�A��Z�'�'ʖ+L�[��H���1Lk:K}��ڻ��lհ��;8X��G.<|��MN��?�BŖ�a��_�.��
�?�n�0oNa�7�F�K�������K�n�YZ{E�d�2���������.�C0�ļϏmw��k����u-#Z]��jc��t�����ʪدq�����#�7-�K���%�`H��ڹ��@| �~���+h<N�����M��Gu>�Na4�q�& A�YN�q��P�e��oG,d�KVo��LG@�� ��$��3�'��=eܖ�����.�ʧ!��cj�F˻̧d�6�&�7��>�����E�#��
�v�'ZvnE:�����&����8q:�Tlo������wÿ����	��8�ɻ�|bOe��3g�K6բ;�1�~��������8�Y������?8�ه��g��.|�?}$E����	(�^K<͚L*ƾ��i����z�*\4wצ?�k2/�43�mo�����5 �a��<Qi�mY1AG����NCۦ+>��:Ѣ j�m���f���~��3�Yhp2d�82h#�U���o�Y�r�W��M4�1~ J�P��WI��.���bhq"�<�+��p��/���#J|$�}��ҙO�k}7��A�Y��y�jȁ����D��#��D�|��a��4 ,�|��Z���hȾ9��ʇ!���Uv�����#�9�F{�}fq:\�ʘ��;0�>���P�����D+��K��(������ǌƩ��7�"��:�
y��"�Y�����h)�b���逶�� /N~��S�G�b�V�ȱ=�^��9�٘f.�<�+�	?��"}2���Q�Du��3��2����_3�3� ;�
����[�W��<1��!�Cż>�ɸwѷH�av���t�!03TB2�e�o��戲�Eɴd �^\C����U�h>UaM���v�|W3%��Feg����#�y���_u��x�g�Ӗy�Y���S	�nN:�J��EI:G �a���#�9���'���,v�g.E��&�����yv�I�����a�މv
i��J���/�o2�N�!W�/�o[m)���Bad�ѓR�Z�(&nK/�y������i���9|��И�c!��ؐ5kc��O��R`�J�1(�p� E���`!OjH�i-��.�P�����	��v;߾K*VJ\k��P���l�����܃�Ԯ)H�3v�s�Akߤ�Ճ�䯺��똋�~a'�gC�B��J�	���I��y�����?�@�����������Z�C�ұ�b �b���Ex�XG�y�/���rɊL�V�^�犏��{�x�QS��C21�&�5d����E�ҏ��l�4�����4�ڵZ]��� �w��� \l���BH�Uޣ���@L"@N!�M�1��P�2�Xb�]=�K�w�D{�ny�_x<l�+rHw�񢮝�Ft���N�Oٴ�ʘSE�k�xI�p�A40�s�tʳV��2r���4�̉�-���v	����R�z�F�q��P���	������|�.6܌�tnRw5���� �jv����lW�$���^c���C��Ltkt� �W���)��b��z��ؠW���SJ�� A�{S�%,N�k����=�Y6��UA���C�}pi/0x��*�~k�%����M�vyA�����w��#�"�7O�H����=A�7�3o��>��*�6�3=���B�����M�$Z��cl�[��z�3�L~�]zÍ®ws�S���c��t�2Tqw��RX�d��%��u�w��j�ՋH��jhշ� ˅{8� �Ԫ4@��'H��q�)�C�c ��J�ְ�<���)l��6�����s�Q�+�@܈��r| ��Ŭ�4��U�g��ɣ���h�4Ήd�+����vmj�<��Q4�?�����}�3lD���C����Km͓g�sR�^(��V8cH5&W��s�sxՔ)apq�
�EH�2Dc�	/��x~�Q��L�'�F�\1�y+l��Tʍ�?�7Lmx[nW�}���:���d�a��rp&gd�0��M%��F+�,�d�c��Q`�����`B��꾩=B��8�z����<|C���T�*ߞ3>�R�,����G��ĸFcxWI(�q���u
�;����)�Q��8����⿻�S�
����nW(�D�ǇA�C:B�K��P��P�����h�]�"6����H3����Ĩ`���@�T?��GD�i��E�A\��%������臺ķ5������]�mH��U�!}o�{�X��k������Ӡ��p�t#�z�c��R�*�l�C�5p_G�	�k��Lt�d9NR��;��`�
nD��	��d������&Ds:�`k|�{�Ƿ a�P���J�0k���0׿<��i\>j��2֔3,΁t��ʫ`R�o3'��G`�t/m7a����gAt/�Vn�=�X�bb�I��	�!����Y�.�����J���\A7��v^G�Q0!m���Q���>]�	�ظg����E�86&f��5\��\g-�gBA=�����ٹ������<�9�x�� �ǽh)����VAs�8��b�=r �;�������^	���n��{!�?:~bY��hZ��+�#�҇����2��!1c��f���w-�>�������;��p�,����iI�x,���k�Ѳ��J��96����#�w���1�< �3�H]Gٚ���d2��ۙ�2�K���_�e�^�������}����bj�A/��pI{��ͮ���Bg<�4E�#�#`�aS�
�(r��e���|}�5���+% { +�p�����{\���d�^E���@a�jy��]�ؓX�⇝$6_&�W��K۠"
��M�B�=#�pP�;�9uz���CR�C�8��w�:�S�G���SR����>��9��u�lm�j�<���xPK��wԼ��Ǧ.��|�Q����W����t'34T8+�C6@w��������cW	�,�M��<j��&��GEQO�a��B�KElR��[�����@M(|�����U�'h�9(e"C���咃CLy��x�$�#p�$땵�J��dI1��	��Y���g���+�������2��+�q��BE��k�X����l������0ħ�l��!k�j]p���j�7m
_�+���Ν��p��k�����6A,���7�����SԲf��n�f�;U�T��a]S����PYʹ���V�	�ޔ1���5�yV�R�kz����U@�I�II��G��'B�α��m'�5�������&�����.�X+kC����Ӆ������P6}C���l����� }a���w7�-��/V�x��Y��00⑊�y��	��֙D�1Jc蒟E�a���*+)�+U�Z�J",6�����v�&� j��h.���#f
������ZÝ�	'42��Z���F���� �+.���HS���ƫ� Ĕ�]B)�,���7��
ݗ�f�{7��1G��NِlcUA:P���Y*���օ�C�PƖ8�a�t��7��7l�p�>�������Ο����%���y�6�� ��x��.������[>��
�ԝ5��u�c+��@�Jv��g�%�s ��ޞ�>�Ĵ�'u����Yϗ�w4��4U=�ӻ��&����1�2�x��l�쵬[�`8�y���k�/SƇ��_�yI �vM��3�[|ӓl>ז<PR����S0�PS�݇��?4�C�jta�ګSsF���"h�Uh.v�P�w�B�{"�� k���X�"��F:���_'���Smf�� Lm�O�XMJ��-�,��)�&5�V�`��I�����%��n۱?����:����5��Q� �>W�P�̩�����7C���hga���/�N~�9����Y ��I=�{�4pz�%oE޲At����p������+������<����U"��r��L�({4��tTv֔8ܶ���^9�Q�z�b�:�$? P�JƠ:u�Ho7���<f� ���xpzX̫�����)C@g��y?z�^���H$Ӛ��j�a���w~���^�Mx�8s�X��i �!��2X<xO��1a_TiknE`�R $�%�6�����egkgi���H�0h�M���V��3��A:�8���ÎI�l �>n5	��N�c5�g��,�x+@$����oTۯ.���zn�Õ��U`�_��Q`����7�gy_��${W�b��"0�B��،���`t��c��#e#<IZZz�]����l���P��)��F�zƺ �B���2�k��9�ɗ\�f��F���LG�D�@��]�Mߏ�H�̴a����c`pr"�'e����h}�$������������P����$�'�q�O�Eao�U3�U���Rھ��U�R*���X��U��_�BĴe����G[����v�U��;%Yd�h{��fA�\:Mo����k��=E�\㛨Ϟ&٤2�x|�f{�!���բ18Iŏ6_�� v�;��+*|�t���#+��Wa@�Er,Kw�GIn�((�y\B���Y���C��L�_k05�u�[ch$�`�!]ha�:f�,��8&^`F�K0���'�S���~r���"Z.���#5�`��M��b_�j!I�����"5�����S5z6�y�x�`��ޢ�6�͊��S������Q@��G��V��dr�=���sk�%��E�~V��E�es�5]ՠ�I�0�g\Хq�9$����da=�~v�ANTX�bv�Aa��ѾeV ��5vr�B����1�������Y�u��Q�lYH� `yd`J5nz�J�����E�f���_�;����g3S����g����vYC��T> ��F�JD�v)�Ϫ�dP0��8�!HA�Xxb��-��
МT����	5Y���wrލ�D��3��Y(v�F�fD�Ŗ����}Ĳw��������[G�GP<|�m�˽3gt�������	#01Fê�!ɹ��
��0��wك(�|�-Bć�T`?0�VB�tE��/��T4 �i�Gw�  0E�nh�e�j4�DiQ@�� O&�vU�� P��{��mD�4v^a�����z��N����Ј�W��q%�;���?�,}ؓo�[����fX�WW*��.��ۥclk@u��G4��������R7顚�*���/�$kI�ذ���'pD��`P3&��PNVQlh	?��W]ë�n}%�5���n�f<�+�D����YE�MUX�ŤU���]��w�AvnX�L����XgvU[Z�d��}���e��hz��F��⯪f���a4�א�]��0 �M���L�?s07SG�t,qɋ,�L%C�Q��e(Ÿg��$|~�	@�ش� vj2��U+�Ļ����!i_*����d;z���# �ߣ���ƒ^ 4��d. �o�okΖǸ��Bq��7{1� ���=�d�(ۅ�j�׍G�#�����~����B��D�㥹�T�PVÍ<?<�Zgd�ֳX��A߈49�F�������t<��s�/�-T��k2�U��d:�#�l@�?�(������\�H"��$��r�_��=��hz����a� AjX_{�X_+�%��gյ�c2�"Fn�x����Ԋ()A�X���P] @F<ʯԡG;%�Jp�7�F(�� ;
�e3�
dgs@{�Ā��lP�r�5��'/(�C�P�EvG��u:��bK�K�Ʃ���f�	������ާ��/Ĥ�`�WU�Q��?� �L�0�;����=)˟a=_�۰�*Э���0d19 eJ�6�F��f_>np����o(h�%)I����M*ve�+�p���j�\�Z9s/�b��_x.^]��2"���
~�)���n��)���Iݽ���]4օ'yF^vɎ'u����ƞxNܮ��79D�6�_���Z8� �F����^��\��䎨�N!�8�xz�k"���FGa��p�p���Dy��ĨVG�G.�h�IKt�%ʑYĥ-)�̈́'ѷ���y���D�#+I��j=,;ibc�C��qPA�Rz@m�w��(A�_�D�à����dFDZ�oe��)��&��Ɗ�6�h��#ˮ��z+���D�ȴ������=l�Ƹ�+�}F�L~��,��O'[�϶K߯�I�}e.�]��$��޼��e���I&��[��?�%��޸���Z&����N&�/#�t�}ܐ�Ҙ�dk3R�㭋s͵����W����)_f�P��F���N�GI��F��aD�����bW+z�`�����ǥ��=��*���H�s�ތ�T��:Ӏz���J�P:��r4�٬=����/m��`�U��T2GM� �i��a�I˄��`$����G'��b���!)<��=�bA�]��m�����*������s@��<��d�k�5-��%S�ߑ�Ia;�f��z8����\�U�g�q(�b�c@W8X� ::��3�c��֌�W��H�J{���C$��i�.������9��tNs�R������Q�v(x�� ���`�E2`I*�6�q�d7�Ed'�KnR����p�B�U}�:����)���gޮ���:�n�����W`�\�f�WKA�D)�~��Z��~oq��e/Eԏ���wVY�o\JuH�!p��':�N�9�g�[�܅\	np8�����hzi�G>ed����P�hh��Yh���3��kZu�W7P�`�kIi�ֆqjG�SA囤��O���R���4���9����,��WD+�Z%���������i[�f��A7�m v6n�.�j��!ӣ��s��eϟ^j�������,�n�}�������k��[v�EL$�c(|lrw`�n��K�`��$iV�Q���-E�27%���cg2�ڰ?��:>���i�T�����D?>`���{�������� &g�bX�6ՖN'�H��7�������_��qS6�F
���ޱ]?-ъ�	mP��Zʻ�{��TN�����C�Az�l7UL�Ψ�T��~��E�4gj���FB��Fq�����`D.'�W?�aV�@���Ga9 �kb�*�|a���x1��O�o��ӬQ���l�}�|%Q�Ib��S	t{��c����ŽW��U�9sj�C�DU�"�̱|�1�Ɓr����\��uY�><U�QL���e�(cߝ�1)��V��@�~x�2oTf�ar�?���m�Lv�(Q$�ҟA	����Z�W�1��ʝ���������/��s�˳�M%	�����i��|0�4��P�q�������/�F���Ϻ#E.���^�=!6/X'����9g�{�?WUӌ��K^�r޻�En<B�}�w�+|e�f��(Bˊ���(\�}ʵ���,��db]wn*��
jB��\C���˜�$��$6�ا����� �>?��;�Q�����<����0������&���>�����p
!;�~��n�O��nΤ��Pa�K���n���sȗ@ѓ�&���4{	�ڇ�%��Ph���$?���L�"�Ne ��M�5�]��Ei�|�'.�0�$�m�p�v姲=�&���^
�ʚJ �n0��[d&� .�=$��8��$<�c�-`*�[�h���6��X�{����Bʺx]�Z�v��\ ZG0�k+n�!��N�R�-�dz��;���|Bc?�z�0��u�������"��6��60g�+J>�)M�E� �!A�e��=�<��F(�ZR�����T�,�C 3��1/BN�8~m����Q�vR�a�w�Ό�T˜N��F�#@li(|W�&{��K�~;�5��yv�i���4�Ҁ?�����UF�|�
t�AL�G�"®����#��,"T���[5�B̵I<ǳ�ޅA�� x�&��1e�WUf3�	�K�� ��眚�$Ό��3�
,�~a�S�=�U��~�'=�8�/�U,�:`Ӗlj՗� �dX���2\,(|���և���46;��`Š���3�(�%�ؤz�V��-�V�������Ɵ�[��,�l>����b��Oz��{N��N�
��;:��&�8�ny�e**+w�b�]�KΪG���+|��h{���z���{v�Ɉ@eo��A�y�HLt@K�:�qt���+q���ͼ̱=�T�u�����{
��ȍhO�x|�m?4n��T��R�t�������I O:9�H_�T=2�-�>��`!Ey�]��/˺)��k��z�IM��K*CKblm@{^���C��b�_h�tM�yB~��
`�b��69��eH9�<5��%Ľ��)��R�^��&��o�����m��-�����v�Ĕ����~B��(�4<Y6�A&����;��A��IW��J�n�fxu�gfITmR=���x_�����o�/�v"!?׌ɏfI�~Ż?�5^�]�g;сa��j��6����p��[p�ֿ��vK��ާ��}�m�f�2����T*o��^�ح˙dX��I>���NychRЪ̢qjlP~E#w��t�*x�H�'���Ok[y���f[ϵ- '/y�/m�$B�������_2N2�];b�+�'S`63)�P|0�%(���lu�M�l�)-�yg{�G6���mz$��r�A�̘,���@�~G.�@� �&�x���/����=O ��ݖ������L��~CY¼���:�����/"?5'�J�eqߜ�=�������H��j�a�
z�'�1 {K(u"�ǉoM
B^�k���Jځ/a��7��"u�d�VW4��ɳ�<�P�%��ב����]��8a��)U�-H�G&�ɔIƿ���[}j��I�R^�1Wy�����/gS�x��S�8����ޚW�--�?�S��+Ґo��%��~; $95�IZ��WfPUj�f.0=X���	l�:ZI'ع���[z��=g�c>Y8aL �s[O� � �y�(�7�&���ag�+��햝�u��PO��kLVRs~����w7~yN0��i��C]E�jE<�06��|���� ��*����hj\f�x/]�\��	���_C��n��J��ف`@3�-�\��2�t��w�Y?�"N �(GoE�֤0�:��Z�/��ڄ��5$Q�]�y��6������a�oo5�)�=�x��`d��N�9w�4�D�c��ŒkQ��5;��~K�w���Af�΃�Q<Bo n�*�(�`� �b�a ����ֶ5��po�6}/Ű7G��J����ݒH��Bc%�
-�I���=06X�h�����?�QT;jO���o�uř+�,�e��
�q�[��3��I6ly6d4�7R�Y��Jx:�Q����pZ6�-���,�������+ւ�Ѧ�O��ְV�>���2�����!���ŵO  ��N~����ě����}��K�Q����b��{@VJ1�#ޱ��Y����wzS�}b�:$m�4"�֯��	r<!~��������x�g�����QO'3e���ع�x��	��j>�ϴܥ9����9�t��
�������U�f��U���ڎP�	}�\�V��4��A"Æ�n��mq�@���0�n�bNo��B�)kK��&�x!}�g^�A����c
+�@։��	�2[Z	
KW�m�a7o������?���O�[�@����@��)�#ɓ���h�(d^�������e�����W��2t�xf�.�>�L}Z;F��x��TPpz�P7�De�8��� Mz�"�bm:%� ��7�(Z�B�L��J�*w��~u�����S 3y&��{g�h���QY2�<��r?�=���u{#A�N�
2�o��$Y�MlAt��-�X�]*U��Cdu�e	��mc�ƺ�?W�+:�#K�H�q�J�1�J�:��S6���p��q�l�G����	���{ 3S��X���	�z��|N��8������^��z��.L�I�@�p��IW�'�����crv�@C�'�"���FQ���fG9�K8��*s��zu�]o��h�ٴ�J��E�	�	Kg%��XE�ǉ�Z��^�po`��"��)gC{��aQ�Qj��c�ݲ̼:��M�ģs�=�u z(�.	x���d})A�:�Q�8�ٔ� A�^-hG߬���5�����)��h���v�z���������{�x�dG��=�l�"����_���_�X�pɢ�!A��F��`���Z;1K��dDe�KaL4&9ί�M��ݎv��cP5jrBsX���_�ëi�O:1&Q�I�\�����u�]�G�M���	N1<��w��[n�%j�j��;j )��W�](zA���FB�ʹx��G�9����o���Q�pt~I���yLL�\V���>��=�=m����O����К%�?�tkK�����ita�ކo�OI�ڃg/��0��\��X"��+�%��}1�L�jY8�,�V�8x`XG4Z>�XjV�
��!O�ġ9Y3_,�^��!���	��p#q~V���b\,�����.<v'�Nm�x��Ie��P�J�#���h=�
�гפ ;�P�ϕ#(��h��guɬ�±sT�d������PR�7<��c�raL
��DJd���
1��a�

_;mߊ�@�QVZd�0Tۥ��V��SVh�t�^8��Y�@��v�qh���p5"����$��D�e���<��G�5Ѩ�D�w3�ꪁ����mA���c#�+h!N�%�*u��'�Hڱ[.d0YBny*EpA���rU^0B�V�Lg���d4��|��r��x��sg��?!��^�Bs,�*?�Īt"�.!~[)=�넓
v7��{v�����Q�H��܊h�
ÔH�/��������)&�ͦ������
Ȑ�����kB�5//��ǲ�2�㽓� �gG���Xd�m��4Þ�@��1q�imGg $���8��Y�򜯖"�ˇ���@F�(^�)$ِW���MbpH��ޏ=�K���8
�]R
N��P���!��4�h:2CZ���\�����%�'V,�r�#2O���=�QH90�	�[t�:A�/]<jD"�կ#����m�!������k1g?�v�ҵj�hɕ``2�����!y�8>	&� ���[�i,��6~�)�ؠmz����H�g���u�NІL��Ջ�q�Z��ڰ8n�HR�!��G�X���m]ݘ���;	B�.�3l��>`a�0�lg��>Ioq��q�1 L����-�P״�v�j*�!h�!]bb�ԎQ36���"������U^.�w��@2U0��A�s�s�'e�2p<)k��+���zr�b�Z�v�d�H{� ��+��9*���D��2�����`�+���/;v��W�/�`H���bH(��<�X�1�L�	I�T��~�S�ޣ�e�T4"�p��0T�A�":��ο�[;�$@Ol��.'�1�M��Ea�>A�.7z����L�ݗ�#�(0�s/M�233tDҫ�4��x���l�=%�cՙ�W�/2�?G�>d9Z�O+.iU��Ӄ���;��W��LDp�S��o�@��z7d������p���ûZ9����ު���N@F$\�D� D�/����E�俾fx�棦)$3w�J~�z�Wq|���7���@�o�~��H��M�B�䅥�1Hd�����G� .X�t���S�7Hx1�t�w�_X�i �ZbA덏y�&-,8{��}20���?�d�-?�tYG�j"l-SYX!2f�kǠ="+�0.�%��LE��V�oV�-��X�8.u�{�y�Yd�jwM(M�Q��{@�C+�~�oJ���.���v(7�B��������4G�,N
)���n~�FzE� m���Z�h�[�X�8�/�kc��s��BT��ű(C�f����}��T8�Q������C��H�2Si7Q��6�5��O������e;�$Y�Eo*��C��K���~S�������I_���>K/�#+s�rZRu<��CQ�wm���sx$�OB{?	��x͇���E�1M�b�j~�>s���s15s�M��ieE���sܟn�R���p��z��C�g),��V��{Ml�x����0�n�0�QJ���w��5�v�k  d$�kM���-) �� �kq\QyyI�.R�5Ф�(�k��s�nW�oUs�nRrS�g��=މ���vѪ��|�
}X��|��!�Nӄ��C�TnZY�H�����:`J{�
�"b^��2"�ˀc��$���תD�e�t�m3�`\�O4P\�̮G�)=d�����x녏>)/ ��n5�CIˤ�t ���?,h4,� ��)����8"�S�+]�?3�u����K*y���X�,8�3샀NKoVC�-�����_UbKO��H���FyN�k�<���F��q�Eh�о[��^ E��{��k���o����ӣ�M�Q�3�Fo�X�B�q��
�?�>���:��H��}�J< ϣ�EW�=�q\ �_&�7*Ӈ*��D����Ͼq��fЮWm�Y�m$�6�zGK�E�����!��ay`<��f!�<D�γ#�[I��v ƞ�'�&�f��kO�w�x��8�u`@l�v'G.C-�6Ӯ�5��D|s��46��ciU�H΄�@���Z��Y���͍$���w���"�"؝���>(�E���TY7\���DSc/�G�#��g=�t�+株��?����[8y4�#�|��T��⍄�8Xw�'�ߗRr$�\Τ���:� @a�i���ܷ���8����4k�I�1�*I��xA�A�j�C\�!�W:s5���M�'{��ʱ�����+��Ձ��z�B�(!S�J�ӎM;���� �+mW�C���!��[�c�`����i7�kU�q�lƚ��QA�$z��sH,�e�{Nɡrjd�K�̾|R�Da� W#�	+��Y�-�
$����*��T��Ԏ7��M�ޒ���f�/���D��w�I�vd^/��~����W^�Z��v%U�7��	���G��sDn���rx
��)�²8�F���<֣�o˥��</��J���]���+S�X#8�~�g�J��g=n�8	��G��Y����ІS0�P!�[.}��u�}�+gqacE�pH|{0	���B,�{UB�_%�K�d�abj�?�>1v�x��>1�u�)�*=�_�T���F�Ǡ\�a3��2̷E4=*��·�T�f�%���{���	���7n���،��|���g��2��9u^0TҘz�G\��@�B�+m�__N-V�睿��<f���Ǡ�@)x�{��|sW�yh���c�'�K�f|eZP���?on�G�5Z��ޢ��{�lJ�ę.2]�(��!��*q��tX.;g�?R"�&���p��Y̕���ӏ�i�~tRE�"ֈ��#��p�c͘yXTf�^��&���5�*�t0��hǠ��>�LA,`����0IxJ0z��?D _G1f޹*��"y���'�3�J]�<[�p�o�L�sT��n��
!�KR���vڿ�bf�}Zf�<\�H�?<L{	�_�ő��7��y��������/�y�jn�=jt�p?g?�v�r
χ=m�X�?��Ǹ�z�2��i����n�}�.:;C���,��_l@�C�0������o��W�ϲ��刵1��x8����܍+�����4b��BD�n�Ջ�L��'xs�yo4�de���kJ9Zq�V��c��#ʯmJe���/��a��Y��s���aߏ9G�sv�д�Xr?ц4�d}|/ݩ��{����B�Tm%:�`)��H�qwOp3d��h��9�������d ��TǨ�R�_���K[J�;O�
L���qn9:Қ)u�n q^bW�Gaů�">�����I�u�ό�1�0����`�M���N0=�W�z�hI(����P� �8��U��AB��D:���u�G:�7O��2CM�5����޼�$g�����XQ$�M~���wtzڶڀ�5��Z%OG}X�����VN�����fi�q�-��8�:����j�J;.!"΋ZsVY��c�掠��X�K���a��^���
O���g[��_S�߼��\{Z9�.����W���)F��� ���T����'��O�ַȜ��[ɕ���W�Z�Bz��C�x�(�[�Gh<�T�u{�.Οc FnT�,L��n:-]>�Z3�����x@�p�n�����sQ��/ju�&C�V<�$]�������gY��>k���^���׾��:�B�����Q����]���>L�W�{��7�{���PV.����Tq4�
������9��r��<Z^M��B:y��  d���`���c#`��?����@Rw�S��6e�P����n0�h� ��ۜ�S��B�I��Z� 	^��|�*�D�Q� ��x�:��ȳ��hr�z�⎊~ak��W�Y:��c����v&�r3Z̩D%��z���z��%�����+C��t��O���@�6�Y5J�R��]@��N"Ͷ^:a��$�����63�4� �|F��t��=:����?�ٟ�d��n9�o�*M�%.�ݧ�	3�����S�H���Nӊe��9��Y�w�9�5�=V+��Nv�U�Ð�Ÿ_v/,V�vl���E�ȏg�V�����8�2��^S`�!���H�y�}A)#j�xj��֜Юht�_"{��j��[C`ךo���oX#�mx�Zr��g�x0�(e�V��� '��̙��X*ڭ�������?@���bTNH����̙���d1�PB��V=���	�?��͖��$*AR'��E�
< �@��@P��TPo����� �2�Pk�,V�&�z�ъ�B��l�6���g�K_Rx)Av�dcpoLVb�_���b�wQ�����iX��nɴ�2��UBK��|�Un��m�.@
�g8T�S�D�����y��0d[��lf�n�?5�wUbp;�#�)�� ��]��s6�ឳ���ƶsH�s���Z�%���c-tb�Ulɠ
@�>�?-a���c (�x||��a���lQ�S���������$����*���}�CHw�^j����PZa��i�s��m�V��4 �S��>Av�E�C��ؾ.Q���Z���02꧊�B��G�0���BT�=�lẖ�l��M�Z�x����������h�"u��{��0��8�2����M��A��cl�<�@��{OF?�$D(N��A@+�����8�e�8}���J�?��&;�*<�9��y/~>7��t�-<gDpfed�7� �h���ì@Tl')��|,�l��.3�Ӗ�\�� �qi��"Nib�&�a��%cY���������◭���l/D?��	����Q�T��9.1F)�ض5AG0��}�����V5�=�)��l��)R(�$]��RT��I�۩����J�'�I� {d������&<�s/�T�4N������lHW��&�!�:�� �Ln�C^�_�5X���%�t�-���> F"��j7-z�#��5?�-�!q�FU��W��Qe��^��$��Q�*d�2���j��\�gI�-w�`#pc�팀�詃�п*Q�zsi�r������r󥏏���C�x��������˙�5�sF�h-� +���1�ա��\jN��NI<�F��&I�q��U�{�|zY�WK�L��n�R�_��t�����6+�U�]t<e�`B*�Y��;�ˤ�Mg.1Z�D�Q�-��re���yn#�U9򒀬b�Aʴ��~��	���ٗ������� ��x��{ύɻA)��ŞH�����@�*{[���_���K�v��ӕ��ӯ���T:%~E�*����d��CL6��[f�`Oj�e�K5M����(M�/��jk�^�H'r4r@*3���?΍q�q�>t�(yA��e���J$�:-�>,��b������w���`k��q��f�������.

��jv�1P��?�H���)/������}R&_��4Z����2�c-�����%��kJ�h���n�DCAP-�;ktPE��{���u,�J��Dj~�i�9�d3Xh�e�^�.���Κ©�B��K�K|��X���Q���鉙��x�ƪ���Z]�j��|w�������HG�q\}r	4oV��x��ݸx�ئ0��WJ������]���GIߗH�ڡl3�_�;F�I\�]��+�d?��_m |�/�r��jW��hN�����q�-�< +�r1�vE�<��ߴ�N^7�Y*o6)v3?H5������1���`��#���+�	��a���E=@࿼byOd]w�wC���|W�j_/��G4��x��~I�W\���B����Q@@�9R	䣀~=3C��Í�l0W��H�|&�������ޙ#�9!�K�F�}�2��f��V�
����aR���v��!�/�JѪ���W��↌;�r��^����'g�eA���[���e;!t^ao5>Y�Dב�q`
>kQ$���3υ4a%墠$��Fy>����vц�JdZ͞
���`G���-��꓾ �=��Y�a����'��)\'r�Xl����Dc�
hh0O4ow����~�8%����P��J�_�k�^mQv���[
���i�͟�������U|�&��T�@�s�d��>����{Gs��6����ÚH���hS�e.1�}���DT�b�B5�5��q��q6�3�"a,C��~�E����C'��>>�V��� ����zB��;�*��ak���/���Jc�}ɵ��߷���7��*jk?����c��c�/����l�b�́_�Y,���#3�+�~@���lˠ�?$�A�O�|�ML����d�+�3�u��	1�? ?�gzw����%�fqx�˝F�;p�vy1F�s�z;*!�b������PQ���c��K�$�9������;e����?��g��@�,LϤ�j�RN5:)�-ϻ�&��.',����u<_�'�d俞 �3�^�K��xg �u��bga�w˼#�+mZ�Xi��{@����tB|�X�y͉a�p���'�n���l�lv5�"q��ˤ��1F��0d%([f����h�KUF����*�c�J�'�!��.)�Z��s!�+@x潪�0;�n�3��V��$R����#:�o%��Ò��4�f�Ĝ�'�*����c�v3����Up���?>!F~��&�� ^[u���a3�#���9;H�chU��BU��x�a���e��L����}b Ճ��U2�}���x���Sqk{��F�`��H���2�_�,M�����:�N�H�#s�75��6�{"_$�� �~d�`�7@r��)^�I��S�>�|���!������b��%UX����}-��=|�14���l��vӦ�4ŀ����m�^q�9���\�a9`9&g��;~^9�~ڡ�FdB`wk�p=ǥ�(����b/��[�����A��ܪ/p��m��y&��p+�t)AY4�(e�D�ƥ�3��1��K��������V�P!N���ěZ��}�{d.�璅�~���!2�A ��k|�+���F6�H�� �4sv�5�h!�����*�Yd�t�ES�",Z�o_��G��<������:P�b0�r9�y�B�������҃��p������M���v��nΓSj`"�5��Qp�2C���+����<A�DX�`uO� ���.�"�����
��Q�������'�I���{Ӫ�[rlaV4��0�ҕLZb��+jm�2���ôG2�u)&� �k�:nU�8v�:vz���Y]2CPT��7
��+�����R�J�6N�"�#"1���$�f��$p}��>���1����t?uj^�T����O��F��>�U,�Z�������C�^V���q�Z����K9���l�(�Nm�n�ƅ:lo����=VвkA���9&z�x�0�`�c�8P��=XE�rUi��io�����%=S��{�� C��W>9 -B[�ћ}z9V|B���6@�X���������1NG{��K��![�+�6N���][)���,35ٗN$ư��;$�2��s*ƿ`�9-���[��/�f�����T�X�j���T�B[!e�J�8��E��~��s�(�o�N:�,�u�z-X5�˪�8x`�N%��Q�I9 ���k�q���/3�Q��p�5.�PC�v�X��iF7�eϽ@X���d�ժ�.�&�@EhLSǫV�Z�?��Y���^#���!ٓj,��S�4n��dƈ�b������ť0-�����)�ϯ�r>Ϭmdڥ,���	�J�IF��+��ƤY�M\�*1tc��̪�A�kD6�(��ʼ�&����N6^5<�Â!4K����H�h-۳M���#�5%�Xp;ZEK6�����>�,����7;�e\˒+>� [p�U��z�[%{fU�[���9'��X<A���%AM
"���U����O�da�7�>��.�[s�=y��`��|B�q��&feyT%�'���;�%�\��iA�l�I�ʟ�[�v(FKc�J�� �d"�br):0�!�8��=�<4U��$��i�m�%�9a���`�O�����ڐ�w���(���:�X��7�H��]hAşpļ�lK�v�1R��?��������{2&���I�[�YX�B�G�m ڃ}��5]h�<�~~5�-�o�G�V�Ci:Ь)�~s��&���,e���[��M�Ej�8��B&�����J�5���a��
(r3�,�l�p�g�1 -��Ag"(��Pâ��"��bb���*�W�>^�3G'�w���ş�\ں��R�]v,qt����[���fH\��؉�]�PRar�y��P� ��%��C��F�D-�A���œ1���YN�9������4�����4���2yQ��q��o\X԰��s��G`ݽ�zf�����Ith�h�0����U����׊�r�bf�%�*0L����w���Vӕ��Y�Dn�1��Y�-:�mN�W�c�α`Е9S&�>�HX�ʹR�J�;K@9�O1`T<�y�!��	�-p����v/ȏ��)�:���X�Fx�fZ5h�[mo���PpX߶�W�	k�n,xV:N���`��}9M68��[Z.�����|�a��w�*Y���.���"s$ ȳ���E�!���ќ����0μ�14�M���L����A�_��B�������@֦�$���]���+��WX/e��a.Q6v��#��7/xф�W�4��粘�о>����17���o���J\c�d�a�ܟC�j�Eg���ŷ>?��SB��@��q��
���('��!t��ǘ�i~R ��E?Q毡(��;@���55���lYI-<�j�ܬs�6ktS�A��TW-����
���
 z4UAL�����)ewѦ�@�t���Aėh������R����G'�l���)j*���E����B4��қyBǹ�Od63�h5@��݄/ڒ&
!�n�yu�̞@K>)�`~O>��҉*�ܭj��']Yw}	L;����%p���_<o~螀v6�{�Zo�S����Z���!ׇQ�|�g�~�H-A��|����r���p���N������R'��&��u�)���L�lu8�	��u q��qF>�2F��P� �F��|�����z*d����,N�Y��-�Q�c*�P9���t���\<���Y��A�5O}�)�����h�͟B���mQU����J�=`�.�v^a����'�'�;̱�oKt���4�6|��<�r���|��U�u�!n ��P�p���&뱣��i7��)��i�-,�J	�X�� 88��Kk�����gz��<[��lFe�����o�{�"EP1�邝w7���Ö%k�����}����b��c�_E#�Y2�#�Ur���,qc���`ع*}|mőJ� �؈i	5�԰�_}��N'���r�t��L��M�v��KE#W @�D[̱�A�C�ݼ��x�(V[�Z��&�P�;z���f$W��sp���K��5�'����x3�C�h�I��2N'%�&b�h�+�+[8)�[� �|����'�i��|�:ڪC8J�g7@����f�v9&�g�d�p IL�>7m�J��"����)N\���='� �}��a�'���������#\ߥw���dP���:#y`7�r���ဈ3�a]��i�Â�Y3M->�r���<��tp7�w�/+�����n�=�2i�3zSb�fG(13�`� �)���j}�r�0<�>g0��7�Խ3�!׫�D�?Gl�u��'�)$fYgU�y:D�z�6�8q���Բ�I��^]��T�}����`ԉc5��pw���Qy"i/�Ti�qN�N��]!4Ϸ݊.�+�En
��Hnx�*I�r53��e�ճr�>7�e ��uz�����>�� �����u���%q�Z�$��L
�H�&�\|@o�4��;���hH���@J�ɱ�L���~��~3�CZ'�5���G��r�c���v5�(hv5����FR��}(,X���g'��mq����	����SeS���7��6Ɖ-���=�3�����I��<�w�D����b��XVd���p�q0���:մ�:����+!�M��9/�g���OZc�k�VU�Ǘ�%۰`{:�8XώF%�}��Z�۴�/����wbv��2Ӹb�r7qz+m�揘�&�rʬ�;����]���@���pnB	Ql��j�ce>��.`��p��[
����3�7|��@���hȦ�����Ƞ��\�u�G58�p゛A]+�|h$&e�ʹH����ȷ3(��8���+�G��a��2���-����U��	N����|O�G�e!����s�}�썒�q�UU"�QX�_�O�}���3p��.�QR׌��PW���>÷�����r.w]?�������6( �MiІ7Dpy��~����7|�-���؛��K�!PeՄ�dƽ� ��� ���~�����ea#�Ktc�9��� ���X6����g.�rWj<��)��
�&��`�k�9J��I@P˸����F��Mw�x����,tU#���֩"j��iA��N8���Hb�-���u}U�M�7���Gݣ�:���4��fS�.q�Aw"�sB?Uִ�*��J>�S;�$��`�Q&�;6�[�Z����oh}r�z�XH��ͣO�����nr�H;�(�:'$9�����bo�6�5Vs#\�Ob;�7�i���=�d"`r��z��%5%~ϖa;o3������>G�-�	'8���]P:�dS�4�<���ʠ�^<ڀ^�J�zP�@ߑ>a��.WGS�=E�Z�hy�j�8�/��K¿���g��Z��j�������`j�� ��|��)|�z����D
-$���R�8�r%�˃�I�5AR�Cl�x���<��p�j�@)-ZA&,k/��Ej���wX�����{�#��e5�@��,�M놗�4��@>��ׂ���"�T7Zuŉ��7�; ��r�7�Iߟ��"�_���{r�!6�$����=�}Ng"JZz7~b0��Y�;�6��e��3U~ĩ/F��ϛ`���_~g����]$��8�]�.�p����Gi��s���X��AfW���)��<��B�ef���0���&qɇ'�=>;L�D�cD��)EG-9��f�S׃��au̿�zx��*�]��=0��ew���kn�ϔ�e!����6"������AXWE�q����'�t�ڑ���Ѡ�H_xQ������ގB��pZd��5�iO�����^�S�/�X��.�fߏ,�hܞ��:5�.kƼ��qԷy�n�&,:����}��+�����ޢ��	ʆV�w�ƈI�K@��r�^4sш���r�R P�_��rL�� ��|}M��P*1���Ѷ�~G������8�D��3�7��kHe��4�������9�'��u��.��"��׫C��8%فЕ�m��gk������D�"|�.mo���0��)M�"<g�ӊHQfXn�gfYJK���U�!�.��|�����ͬ�)��g4벸L�5���_F���`/5����'ص�w���̦VJ��IT��l���Y_�φDW0�\"�"�v�X�H�p�5]����=�,l�P�f��ۮ�m�P��;p��W�LZ eu���>�+��+�}Om�dO ��!�2�D`���7yC�O����5m�G��F�=�����j]\��ӯ������n�T�Ȩ݀�Iu���Vt�1^; ��E"���5�?��Z���]�7�I��C��c���߫��4��6�/fH/	�H��ESθ�m;�.�׃o.%MF�9��Q��!i'�ڪ����g�Nh'F��U�T�z�՚.8���V��=�=jiԟZʬ�^M���>���&յ.��RÚ��yX��$�jnױ�#����i"��;����52�#F����������u��dh��FG���1%��%��UhL�/v�٩�sLʧc���j���ܫ� �x�w�����]�|7^2m�aP?�@������ƕ��?�]k�B�;�&�빽G&�$���b�Đ�P�N�0Za�q��FU�d!ݞ��VXo��mF�=ײ���ܭο.+N�ʴ�6��g,���x�㼷L���,5y��'?k���o�|��.��F2K�b�I<�Gf�n�H��i��R�*�q�:5w?�b$-"r�PG�䥹zާ�9����=�����m����՜~�CŚy|Ύ���D���T��)+Ŷ�]0a��ZQ'9d~����M���0���<��cr��}el�G��ps� �C�����&'�v�N���,2wv��g��pT
���·��sh邈K�na��k�ݶ�o�Bq�^�����(���K�r�6@���u�#�TO$[Ɋ�t��l�R?6%�+9��d`�aU%蟝�R���?�ʖ�9��\5ŧΟ��9����j��^8e�jӊ�S2��'��u��D���$�1wj��K���V:�D�T�&�Nŭ(N�Ay���ʝ������u	�Q`#Q9��X�S�C ���JD�?2���3�	��]���,�2o)�m�G�����\�F�1�:
����b�4�5D�,+K�2�b�T��βf��nR��5��b��33Kg�ǵIU���g��]n`c�J�[�2���~��a�`��ƎuX޽��lD��m��@)&��QhTR#���z~���F��4T��q�q���r����]?OP-�Mt��)Cղ�D�#�"6�1�ޞ�=���R��y�Q���f0��i�R�t����q�|��� 9�Z����[��ƑU7��o��[J:����z�^����Ճ)(oܑ$�]g� "d�٧���ҕ��ZT�v�y)]1���g\�L1׼QĀAv=��m�Xj����<s�F*�7�ޜv<�@_0��(�-xd�<�8�%�3�`��Q�q�UU��+�w׷`�t4ُ!+�%xI��C����rF���,4���SF(�OqyA!\���g�]�7���KF��A���E�>�'NDo?�&m���t<�Ƚ3V�QM�h4�0�ˎ��#�7i��10��q�R����\�,F�R���UGҥ����N[nNY�:����5y�EF��v8�Fv�wW�Ms�j���X9*͢	�a�����3j�ݯ��{�(	Ʋyɿ��eϕ霻U	��J�����V稫�-m���i�� &{�����j�ɒO��!�C�Ɲj�"`�����'�d�5}M�pa�:��P3ȠA��.�c
�@�7����P��J�}�<5�M�ڤ:j�x�i��¼�2�����'�#*	�:&,Y�>���rzꦺ�վ�U�?��j�M���|��⾾:�����MT���q@���;U$a�je.SZ���5���@9�� �ч�n.b�e��j��mz/�@��X];Ph�x�R�*�-QāLd�����;HT�����`u'�P��k9i\�?_T���B���}B(�sR�)Cyi�?�ȣM�����r�����T&Q��������w��s\���.37h�J��GX�\Qe�v��r�)Y���=�S�5�>��,�K|9O�To�%�֥��'�:�ZZF��Qi�v�mT}���3l��C�փջ���l,�y��p��;����P6j.���1__a��QX�H:��e`�n@��C��:޿.OZu�i͛����� ��p�m�����&1��M-0��}���%�X�v��A�h[��8��=�4[$ʆ<��R���14m��X�W���ǈ�Q�i>�]�QBl����܌�/j4���r�!i��l���-R.�4~�$I5\,B���"��hV7Vʇ�9P���qw�s����m�L^� .���}�׮er�8̊A��G�������S���O���S��JݧXI�οpxM�˷�7pPQp�O��a���
��Z�1�ީ{d��q���2Kaއ�G�� d��G[�k���쯵,�����֧[k� X�\���rNG��0�� '
�L��\!84�P�8?~�*���ع�,��R�S[Z̪T���fȇk97�r�mH��a�@�Hi�[�{>U��1�2|��.(�s�M,�r<;�x�yW�-$���]�����:��kJ@�1�=3%Æ�CҔ�ɶ�Rr�_r�Z��jκPZBg4����`�2i��`���0G vus����_si'�O@f�� o��b��r�� �Ȕ2�x�2��d{���">���rc��('�2�D��1	���hY�ό�n���~r�<��$�9�x`��]ъ�*�&h��P�}������n hԊxiM�‬�nB��=�8�]�j�{���Zذ֩0+�$\�5�G��J����8"?hSf�OMrGT^� F�m�M�w�J�_�J�p-�'��������܁��\1�$����h$��f]c��Pk�V��r���xR����ay�T\�ӣ�-��M����c]����犢�W�z����2աt\Ӻ�_��0|Ӈ�[���Xƅ��D �C������lQ�<7?�.��>�n�Ra�K��'�s��E��@u4N<@j�M�=ծ��$/�8�ײƎ�H�uNI�z%�����X�E>��"_z���IHB�WAWϒc��@ٳ6��h���t!_�RAS����?�{���
r�>����H�`������l����\T�)�g�2k����i�6�~,M�M͒&&�-��+f"ĐZ����`���liM0��i���
I&���jr����ܳ��d2��+�Qi�I�?�2P���T�5�����P�	��]ʆ�5���cĈC-[�y��0��"m��9zq���8���l���q��?	�K�+���B������R��������y'���r\���4;�Yw{́��Χ��fe�N&�ض�n��"����e#����l�;	�$�w<3ce]�Wl1t�񟇓��
BJï�*,��A�Ӓ�h/jA���k@SN���l��*Ǜ�n6���^^���><�t��?a�<���b�,|���*��ۇ��}��f��6�Q�Ĳ6pM�nl1�t��Ή�Q_S=�6�L9& ���lM���l�:��^X�|��U��˸��F/�%
�y��)m�iR��}�x�P�w��:K�-�]\�Ҫ_N6�����=�o��,�~cD����-�MU�ceZ9%��x�D��&�M�8ޟ�=��(��kރ�*�Ʉ�*�R��1\�\����d#{������>��8^&C۽g�Z�]�p{m#�vyi؜������@�r�n�O;�!�:)���N���l�XJ��p\�L� Fyͮ�o��#= �=.FR7��kMCv�9u�0�=X�z����	,����G�>�ϙ����/B�x��1����߯��c9���á�8��c�2��ee��sW5�J�Ưj��I_ܼCKk�e��Ֆ��\)�7v��}��%�B�;P�������.w��"=��O���rjW�Ɛ����9�a�dN7o�!)�3&r���f���_���B?%��b ��N��j�^�÷˟�F[#��a�Mw��Nj��$gZ�0 ���݃���iG�����틅����<�z�J�((��$��Ά�S�_��#"�sh@"�>��!?�ơ�V�C1	߁���:~w{]>E�G38�%��Q�����Nrb�U�^U�	�q~�m�i~17��\!���GM �����Q�ޚ�YltO����!͇�q1{�����U�6�O=gM��/i�U,}��]�bCdZ�5^O�p�4���p��Hp����î���0�������I�����WТk@��q�y�~�+�nR*�L�g�'�I��0h���B�R`�r�9�t��(���ij^�>��q$y_��>C?
1�!��a�0 ��{3��&�tX��9����WG�d�\��m�8�
D��.��ve����2� �1(��vZM�}d��<D��e�8){�.����5���Ue�[||��qJ�8Lm>��Pǧ�1>s�C�Rf�al%:g���[��z�m]g
�Q�V-ъ\�F�m�����?T��ԅ��p|��]�E�����������:W�u��T����H�_n,�9H�����0����<Wer���I�>g���"ɠ�=���
^��Cy����^����FOt�C_C�ӗ&)@I.:������ؐ�4z/�{p)'>r��@����/l�a�PD��h~/1,g�ć���x���2��푯kD��`X����MTe�J�D
C>���,@�)/A��������`�w�Vzݽ�0��/���[ؖ�|�7��əⲆ
aB�5,���C���4f<fp'��_V2Ԓr{Ýz}���˘"<b��-�y,Rii^3-F�s��/s�~��!xU�;���!=�2O���-JBϿ�&$���5;ʥ�-�mG@/�c ]�S����:E$N��j$������A��T�){j'��n�h �F [yJ�쎟h0�j�Å���ɕ^��&6N�/@��#�B
O�)�	���I���B�0# ��IO�xf����
U�x����^̷�r؝V��"��r�'�lMɖ]��U:`���S�����g�J�(������ �,T�<H���NK��G�$�6b�R��s��+Q2`�PN��zy6)��3R�R/l��y!��#���?�P*���t"{�,G?腌�"Q��/�+���
�iu4g���<УI^��7B�:\	U
�����z�+@��t
�]��j$Q�$����&�\Z�t�C��#H���4�(�9�~[���$�^��>c�])�X�iMe������m"jh����
k�;R�2O�&O����#~�ǭ�tDz�$�PUd��j��~��@�_��VM	�R�&��)$Kh9��F�U+���6�(�Y��J�����d���j,(oP�~'1V|���A �ZG��])�<%�+�][��X�ф?����ѓ��|��S�N}'��!ɪ��|*��>�O�E&;��x��-���t._{�+4ͼ��?�$
I�N�#͎7�:�ժ-�e�Ҙ34d�Zl~�G,���@b�85�Zh$x��,+�#!��[���t!�$�υ@)������ҽt�D���̠��={Ƅo�[����H�jXBE@����ˡ�qѡR{�V�]�γTȀV�2�٪��y�9�Y��a^/�88_ֽ�zl�|kf����U�QA�Or$"OJu�j��� ̰�'@��O�-��ce��k]Q����T-߆o)����F�=uG�H��}KGn��b�W�9�ݙ�����.�A�g��xV���:�qK��ko7�p7�A���&:�]�*"G�ыsFB��v��:�O �K�6D��4~����Gzga�Cs�u�a�!�$w160���g
���ȧ�"U�j��4�x,Ý�~��|�EM%��IY�4��i]��X�b�����D�^�h���R��,�hq~]ė�eP)�i��.F5��gR��2X�;���ܩ�X���;=�vhZ�M���P����!�[2��=�PU��L=�w-?}��[��S0-TJqEy��E�ߜ���ai9���))5�5e3��JǪ���BI�/FT�L�!߿�6��']��0���7Ԭ�� ^.���n�@!i6Y�礟V�&�w�B�Ow�J�{u����9
�Q"Yv
a���	૶X$�x�L@���ew�D��"=F�#�V�.i�(ܽ��ɻ�HV�W��i>DFxKIp��@e�9��sW0��[d���E��l�xK(v@�U�h�iF]�ʶ����������<��Cu��A�B��iҧ����H݄�	��j�A�y��v���yZm��(���mS����U/�tn"�%?��z���|��	��	��k��WL�ᦎ�o���NT
&�
���ʸ���FP��Et7B�Zc�̽���)b�� �)�ʶ\����&֚;��{A�^$A�Wۈ1�T�>dC�c�#s �r���#�Io��̏Y�t�jxԅ=��a��w8�Mp���Q�C���Xg���;�y?.H�܂�r������*ʀo�"�c�v�L�yq�u%�QY�*8�"25b���c�ե�m�'�5�]�PMn�	���L���z1�"���N��)���+���K��/�e\���o�
$�bT�
�6��T�'�R�Ukϟ�N������׵��l�m�L͙�OU�>�|���8F�}�^���۞���8��A/�� T��6���5G�́:�l>��{4����䴤������h�k-���te�U������՝.L܂��=����"��Ć���s%t�T˵=�C1�R`��%e� �F7�y �|�IF�g �Y#�T��oN�F`�	�o���{ŭ���	�iN�Ml�FA"����9����I?��� �7tʃ~�u��/ �"�IM\p#��q41��QE�Oy�1F���_�,����D?~2�ݘ�����]z��ޅ�5�����a�|�&P̫8t�nA�NWǰڂ�	+�	��0��b�:��}�26��<�����uj�i�g�~.�C�g�������O_�d�*��l���HH�=�N��G"�����R��u��N<���'�#���a(S>&M@S{�m�����}���J*�_HŢ=�->��Q;��L��+d]�!��ob1]- ��J�&IŖA3����uv?:Y�Gт
��[KW���Ho��O8"<K�2���m��Ֆ����p�`ԧO�c��VS<��R9�A�t���g�����Y��7|5L�^M��xOu���3�vɴ��1]��I�5I�O��'��+ך8��^�-��q�t��5�ϙo�u#z�a�o�/���NQF$�}5;��x���Sߴ$Z��s���({@��c�Q_����/V%<�׌aZ�*g
���i��A���ėT�,���[��9�'���Y'?j�?��`�f�Z9���3z�p�EM 2�<�~ա��.�S�?����	�ߖK:�p������e%�����n6���w�oۥ{�4B�ew#��&�ݯ �#��%����9�M)ϗ�FT@���� ��14�����_�Kţ�p|-�v�*�Z�uհp��o�Ji�yè68sN��J�aZ��~<�2���V�ZP��+���y��}��`ɘ�L�IrRi@%�HZZ�UR\������C�*�0(J+w��[�JQMf����e�$��k�R��h[� �D`�뚟Kb��Kn��.�[�@���O6��H��)y���}}��P�%�hK����/9��\�BO���b�P����}�NEۜ�ъ�BeI�6��5�Z�Y ��I�zf�:��0��q��ǿ�F�i%Q����dGB���1qfq^��D�t������#�sgn�洰1���Q{Խ�HRO�v389����&�*��^�r��ړ�(�7����'��;a�����+�w#�`�W3����v�|c.W���b�#�}�载�~݃_گ����BB��`l�_��%����l��Q��GC��p�g���!R�WZ*ѳdb�s)�̖V�\�s�8�Ӝ����B^|j�?~�z�Vow���<�ƒ����a5�� ��Z�umF������Kw�Q���3���	[�Z��5�������8��y_nM4d��4����I�K{k�QAW������*��2��I�WH<�����n������@����*3T4���5��>�sl�KK	3��������(�����K�(\\+�����e?~�\ �[�ǧjsϨ�(�,Gz?�/\_:P��2�	�׎������,dM���W�^��"�͂�{CNēK�V>��q>Z�#��8�6P��"�G�%��.�\��50ۂd({b��J�i����Č)f�����v��7�#��_�?hf]��wV�Y���|�D�;�@�S���y).�  bF����޼��K��s��Z��X����dI�Kq�D4�j��>���3�� �Ч4��n}C�O�#�la;K9�a�r��?�K.�Cɲ��{Y�"4�A
��Q�?IŴ'�S�:+���?��\�s��<d`m.���e�����(j��di��dg���m�R�D7���(���i�m9�ay��ve��0��$���9��6̅$�a��YR�V���I�+ʿ=r�+�Q=��l�������R���"��H��
A�H�"�]��vS)S�y%�S����m���1��~T_@R���}͋[�X׌L?=6$]��Ɵw�	�/�O]����<��v<�TyQ,��c���4u��8i�_W'�s]-����j�b��б��7����-���=\�dt����A�?�\��jn�h�ۑc�6����ޅ��]@O n�0�4�{2�@XĲ�~�j}�9��^4�JQ$���z�Ԥ��+à�3�lL{s���5-l���oPk��ރ� �Sv�!��R��#
�GȬߛN>��+$�6`@�1��K����h�L}k��c��?vdkP�a�*rg�p[�AC�	;,&o2��}�;�K�:�����j�(�T����O4�@�h���� �_pl�V̳0��5$�&����Q�.�����;�rA�Ơ%�u_P�`����6�x �H*9�i��O:IU��w���V�p�G�,���(D,Y��-JCu+	���H���V��!�-�����,�s�܊ y;'$4��A�;��`Dl����W�VT��6J�a�Q�8}��2K��h�(`��՞O�w���崢aGړ�z.�c��PZ��p�Eʲ��>D�J���%Ã,��?u��0���W�@���dQ��q}����5�ZE���4<m멸���o��a�ʖ��'��a�Dx=�� �U��w�(	p"j}yB�!�N�[�;�9 �����]�'��wL���6����OG��������S�,If�cjFrDV	;u���fh#�Ɲ�޼���
c\V����"q�C�T���j&����}>Q��ɍ�̔�x����� 2g+�[��z 6����$�}�r����� �|Y1�g]�}�Gl/���t�_$��1E��,�������TH�Ⱥ�{]������1�2�~a�c7�C�Z���ё�r���r��"�*<�� ��?9WJY�ٗ�^&^z�������s�Ls`�+�%�F���V9[��1����4r=�����9cJ�Ӡp�N�4Ľ��(��3�ˤ�*Ov(���������g1��^q�5���]:�t�(��)�B�`ʿ|��3�<��W��@^��s6�nΗ&�p�!Y��p�O�ql��.��
����5r�79K�A��p3b�kK}̳�<-s{WI+�)��7?Wػ잀{[��&����%��p���؄�Wg�z�D������qD�<(Ş�e�d}A���A�~Z�J���ϱ������Az����pa+�Gp<�����qe���&�wӳ�'C���?7���a9���k��j�}sv�}�U*f_�-�<������)�r��L �ҽ�ٻP�r�yU���S���r{����o0\nh��՚��M,'�"�cr3��`�w�ch�fy���2�	��i �xɕK�o�p�ia��,W�.��if1]�a�2Y\���.5|�]m�`6X��*����[Ʋ�c�^���g@>�U�܈oS��V��BT`kom'�	�R�}��7̍j�]�q�6���oM�Ã��é\7�߃s�IՆ����9)}��$�³���?�|���lˍj#JyJ&6w'��(v�����)��;K��YV�'H̨β�Zg���z������eVl��-�<.���Y �E5���Њ�0�<Y^Ň/=��=�J�0���l����1l�k#fwl"�$b��#<����@��/� �c��1 d�z��~���9�::9�~���^�6�.��1�#y�vQ���B��T`Zg�#*�!�=���b������A�+��㱈�%0�_|�%����VoF�y��K�~�Kb��D��3�/�K��״Vq��� (jWP���5��Qq�%�h��7tt���G����ӥ-T���u������'�M඄�D	���t�s�}/;�C:ֹ�`}{�vc��^no��3M:lC�: ��Pdc�b���F?Mg���,{����r�%�Ť�)����F62��E?+L[}O�{ߤK[��xnP�!�["�>
3��s׈���ou~�$"�0��lvH��yH��r8���n�P�v��G��N�P�Ű���7�i�iXn�w��ur;ߘ(�yj���,�¹�ޡ���"a�:n�w⸫�M�zJc��:��թ�W�d��#oѨ��I��%Z�+��i���+�U�=���1}!$:��e�������ȓ��p�78�hb�sEG.t{D� ��^0�~��Y��t�Ԡ���*[�����jz.���a�@�/�*O��y�.��<rR������Y��h��	�g��y�&D������W�������c��e��-�4��%\p�F�[H��TլT=%M�N��\���l��p�eǨ�o�HL8�'w�sO�;�w1���I;���)���'��+�Ԡ2�1�1�պ�&�ٸ��#*F�����D�lR�����sD��{:��_���ѿ������u�f��hf4e2�e��g��׬��|z"Y	!)M/'����=��C���"x骍�쇏!�T���� ���i��'M��gɈ�}I�pJRpx�]5x����>��5�&?T:�A]���>���/Փ����=d%TOQ�I�Ĕ�ξxm[�����[0�M$�cl[����]��E���/ߤ`���yB��'.�L̃��'
�m��d�7��Zn� �:"؂O����Gz=�lZ]>��W�&:�xn-�'Rc᳖כ���p7M'~�Übl��/A���d?�U5y�0����d�ǥ۽$� ɫ��B{͕����g�,��4@?��e��ӈ*֙r;��9"���*�)���*����[R#Vl���w7��5C�&��Y�f�H<	"��'�ֆ1��^�N�{��N)���R�ϑNm4`a������d(`͞��"�S�\�G�s�Sҙ�;+S��U���v+�/�t�"8̅H�o+���9tlV�Ȣش&U:<{8d���"-+�4��`|P����4_
U@Z0W���+��@��j�2I�a+ɷ-})Vfjה���kݩ}��+y��7���7}���n��F&�)T��Hk%�V����sc>���Q���H:���!�����y5]����*.�r�����A�[�|׼�յ-T"	伋��}{(�;L�P	�oi$�	��&������*��%HWs*�:^��^�d�L��'����mO�����p�Wq�꿧�����q'��uf�kx�`�Y~�`��F��0�4�q���b�v��E ��*4HŇ�d8NE�H:�e�����|9�\�B�8���[h�	�>Ӊ�j_8Ý�����_��UiN�v�"���|�~����ʋ.�>����N)2'b����n�{%	o�pcQru����a�#v�p)����re�B�����1�R�md�}#��?g;2�S��ڲ\Ok1\Qe�i'����m]�-st`�lxKǳ���t��w^ Z����?��V����+0�jVLY��@N��^Զ�K;'�w]�E�x�� ���K�ҹ}d��
U}U�;�w���(ȱ�2��ɦ�xz54@V��0׈�wPF�e�+r(ӿ>�[?j�;���F]DJ�)KJޗ��)K���
Ȑ}�z,b���a�2�κ��,)1i��/`�&�i��f���&q�7��x�"/cK�	QܼOIBL��xd��o�?3v���h)�-Q����O3��kn�u�o�i�D��e P+$_�a�����Kj�~N(��!���i�n��wî8���DLg�0��nN��1��s9[��5E��j��h��(�el�g|��BZe�N��L�$zBť��S!=%�}U��>x�T�ם��K����=��GRܦ�)�W[+L���P,P:!���v���D?0-I���rt��)ƚĄs��M���aÞS��i�.�g�
ѵ�����5��U�lh26pACu�,�]�^�Oˈ���;mů��\�o�,����)j�n`xo�(n@�o�Iz|̣�+4�>��2�j��>�R��M�����q��0[�r� o�bl�˛NR ���7�˘8��G�Nw��\.�q&j�sq�D�*��L�<���gD4o�$iH���=��J5{�	QhA�m��Dd6�p|y\���,
�uc�(��rz;Jӣ���*�1�[��m�]aag��1��vfUKWgT�p��3���g���~�b�[�$�� V85ݥ/�ԶXx"|�((�-��F��E0�|ڄL."�%���F̝O��{g�D;�!��7���[��YV�>Mz,j�@�IpG���{ ���A_��iw谑�z���px���a� �c�����{�_�h�q7�LX$�T�C/^��N���?���-;���4t�Q�����p�y|݊���E�'�(�6�}��pUUB��v~����$n6_�>��!oz�LN|�Q�_�}U������U�+O\��h`j��2����y~*��y��/�ԉ��'w� Em��^4�e�?�nAj�� ��X��Z$�yV����[�h呑f8<���ߏ�5������p��/��'S<U��坨3+k)G�`u��³�r	���)C)N��2Q���
z�,
�/#��jK���G���1�sA-�G4|�=�-��)R8�%o�p��^�qGU�f���dS��PoB�X�nÖ�f�"m|%K��l����!�/
W�!�ʟ+�Ο�:�k�j��F[���l���~fcl��Y@���ꝵ�B,�]���{A�o�Z�:���vO�@����@EV�n�)՗��m,ܾD8J��+�	�q�"���_�j�ȞP?�o�m���E�r�P+��_�h�W:EB����˘����|,d��Fs��1$�`]'I�A������ݒr[w,G-V#������(Lu��N���~���¼�sF�=�Z3^_�:[���?yO��}�,�#��j���
t
M�0w��F*�?`�.�F�n�AmlDDB��@_I�Y�/���ڞ�݊H�QB7k��G���N���%>�?����U�"[N$Lk��pک\�����>/����]qҗ�J�yw������z6D�{
CoIG��d��Uꝇy㲧8�z��R�T��&��9$���P�%
s_<����xs�Z����Çz�q��;��IA�FD�i�wt��W�0�U��'�a�I�=OX&O��5�Q�K�Ѯ#��iݕB�n�ü����ﱪ�~1��o�!bK��m�+6�%\��XוM��x�����3ȣ�fݿ�}�ٓ�b�,唀$�ɯ'���-�@���$[w`H�[�
��+7�&B_n	��}���3krQ2j����q�fx� <�:	NRB��H1���7���?VnA��#����-�H��g\�F���8�&n�mg�]N���(��$6D֋���r�KZ/�4�X�?��UU�v�r���z/�y��E/D͸ꬃ堊�:��J`@��b҉�����Pp�t��%�m%āJY�,��[j@5�4'�ס��9���<CwXt��MQ	�Vo�)���P�`��UV�rg�0xl��Q��!hUå[~{��!�h�/5kfkH�X�h�T��y=�v���c-Nk�ҡ�pxG-�����v �I�_י"���<�&����Fp�G6��'��f�o�]��x�<Dr��u�S@כ��)JDe�8��7E��<x�g 0��'��7�G�gy�!�h��T�^�"��ìr@>8Ӈ�ϙ�CH�[x�������12=}O�'4��2�cH?�͝Ͽ}��4�S.%�V]��ɵb$�?���)�]�.���Rr��eth��p�P�A�Z5����jm�>��	GM�EU"vE�v��Z��w-�sv��
����3�������7^!v�U#A0�Ј�r�����5E��7-�2�,�î��wu�u�����]���a�A|��`�ƇL��bް� �T9�a���ɢ>��eGN�GSv�`P�h�'Z\JIs��i-��:7��� UP�o#?���
7��'�J,c�t~(T#�|u����q�|l�q	G��Qbk�=a����O}�f��֭-�����iш}"���Ƒ��lE�|3 !�����l���߄V����=�W!,��~(��c⌭����"�0�-x���UW�6�iz��'�n�0�J�W3��qJQ0vdޟ�> \�)d��/�����r��V�֊/���/��pb�7��o�(��Y}��h� ?#gP/\�;XUI$�X�p�j��)l7�QR	Ʊ[���������M�� �3w�,Y%�p+�Ǽ�����HY���U��Ric�,��JH���'ֵ�Ls��4jQ`{�N��Pm�G/,�6�~������e��#�@A<��j�/K!��	�L���O>ޢ�07 ��G�pH��тk�(�ڡu������b��%����j���,ZQ;�ϒ�S�ɜ�8�iW�җ]De���>�P����d�]���Oյ��߳W���xA{
�`o�\7�n�3�G�����7�:�����6&r��:0�3.�	���s1�s
���߬���!�qw#����ix��#s�g^��	C��ԡ=��5Y~��1�fL��$3�D"���?qӗXA0[Q�b��^�≋p�;6;ʉ�]պ��7�x����&�@�:^�ת��������|�S�Ǧ,ˢ��e�@����ϾUp�������۸����s����G� w4u{s��p�¼��/"�"y;�m�sR�HK��V�����ڏ	�9��ó�r�)跁�#0���ג�Y�o���������>j]�_Q~�w��IT��.r���'{I��'&�*�ɛ�̡WA;b	o�1�]I����
L۝/���4"��|��NV��N�����yߓ���Z�lð.~���Y��H�uyc�����]����9�b���w5u`�?�h�W���SH�v��Vo�(]� �v�<;Ϙ�������P�����,
�6�i���h6�:�����G�r��oo�@H�� �:e��J0HT�m��Kz\!vԨ��!(�b��Rj������]�b\Z�	��ۺ+�[>��K�����e���a�1����jjG�j(`�[�|�t�Ҡ�x�!�J�X�����>>Z0jL����XG�aӞ@��]I�zP��v��(��/�d���m;_9]g�Ư��3�Z\�`�urj���9(��7�^9���;5E�p������vhq�V��X��v��
R�CO(��-g��pUT����8���L�1}	SdP'R|��v4o����O���U�D�ꚭ�;�k-큆td��y@F�ߎ��`��t�W�b��2?��*:����©��!Tw#�AxK�FA���]@�t���dWf�%�8�R0(�w�n�~&<�~a�slr<�^�ɤK��/ړ���O(�~C�oED5u�'r<�E���muH��8q�`�x��e>�u��� ��t�2%w5x&s���B��m�n$��_C�0�Z���<^�a,�6��i<�`]�wM�V����u��t�ڥ�ڣ_��3��.8��*y �0މ�X�X����F�]�5$xv��W+���@���*}�}ҥ����P�s���!�/0�J�˾�����L��j޷��#��q���Q|��i�[�Ŕ��-)��i��9��K�Rj����ڝk̢>;a	L�8�(��TOq���}�l��"q���>��"H�Ԟ�o��#�a���]z=܃��|ߦ2a��?rv�,�*�H�A��k�"��pH�ӄ���n���B�9����4S�w/��p���vz�4K�\�H�E���0!T��њ��,^t�L�/�B�gX�S�]�`�����;7.�`;�Dz����ъ�i9g��gI��1���[�m�ȧ���e������'�\(��J`���QB�s��N|>v�9VQ�̤|��Z�K�|~�O2��V�y&|�8�&�Ay����~�ƾb����_M�7Te�zWl+���fr�Z��$��;�")��T����O0(���B��eI�QUhUH']�.lB�/7��-�"�ۢf-+�S�֏���Nю21�u�es&�k�<3k{��U�z�q���"M��_B�6:�����z0�])V�����̈́Kۭ5O����?�MbF�K�kު)�t�w��{��@M���0�� !�����c}�|�:�mP�>B�f�zXν��/vT��]����.������&^�g���ѱ����>ǁ�%/�~�({��B0�.�$ͣ\�iaS��7��r󉋼0đRW�~���&�>�����ք��[E�2�h�q
��Yg�2��꣡¿&{�d�����8��Lˤ������l�j` C�lM�͡��G�b����L�EO1�P�4)R*3a1ol~�JH�HG�e�V_�4PC�(�[�O����fƑ�8��J��4�N�,��0� ���P4������ Nk,꩓�\�ꧢ}	��}�����xk�֏�'��8����e��T����9Յ���Lu���5����"����2q\s:��촾4J�Ey�����_�0`\��_L�	�K5-�Z>��wJ
�lwO��匦���!r��H'�k)jv��m�{t��	�|�g������f��� ��74�3c�?����X1���.n�|9��dm3������= �`<�`����Y�U	��.�gJ4@�񕌺wdj���ʘ�j͑
D;(� 4�x7i���Y?YCG)$��'�4�6��H�"�����2�oQ�T�s˼���a�j�I�MN��y���g�o,�w��	6�ߟ�x��r�ҹ�2Z�0��� �_M�����j�P��2��?q֔-�H�8����9bA=Pcf@�j��{�P;C�I;~wRQ�C���c�WIܸ�˾�{���0�2��ݤ"�O����gw�hl��n��O��� '�V�����q,SJ �τD�� ZSȜGC69V�Z%�f�^�L�����r�P�n|���k*eM/��Ԁ.���.�\�5��Ot��
ܖ|T6�nĆr'"$���|�q<0���LVxu�b�Y��\b���_G�|]�d3��<���90��bU�rZ�QP�F���Q��&��"�I��u5�h���	��Q�P�Y�H�K��� /#�`3�r�L)$�E�c�ha��6���W��[��P���rc��4{�e�s��#Y�e&�q�,�����k��"ͦ��%��D��Z�Б�wVK��DBQ��E.:V7��J7�*zq?k�����ERp5t��Ű�o��k���M�w����t<��Y��e!�ul+7�i���gu��:�:�Nt1�"t[g�!U0�q�Q{�y3Q���|��o�g �{��wت*��S�g��ͭiC��ݚ�f����mk��l=tt�����7�3�)����Q��򯝐Ҽ-�FcĄekM$u�&�J�b�X����7���O����#�sr��~��n��D�y00���qZz�7p֜ྫ� ��f|�F�������Y0�FD5�	�@>�ϸ���Г)��qS:�o�]	JU3@tdU��P�vڨXp�O8�%?њ��w �z�:��SEp�~q���{^j,�*��n�������t����مu_�������!0��yԉl#��T��m�R�� ��K��C���~
�M7M@1����!��.i�yy��*Ӎ�� �`]���7����§@�Z���l=G��V���s8
����y�p�
��9Ω��1��!#�X�B�n�ZBs����H����� \����JTW9u)�(^l��1V�,�~>%yhH|H���t�w���q�����8����D5G��p�nWE�.Y�+Y�6~_=���g��9CC&Vʼb8�`=wZw?��-$C�%[�cXŅ���鋖�<�&1��Ն�s8Jgq�r��T�)_0���r��=��Zx���H�,K�d�9�@|�Am�G��K���n����˳(]�]Nm��eZ�q��� [&���J`E�?�!�ɼo:��m�"�����)�	(R�~-3����`��@:1gXpNFӀ=��5�����l�!O�g%Y�(Y�� �H���z�W���Q�����_��Q�\�Nf�@�����5�* UBt�VP	V
�ӈε����\��l'R�B���װ0,��	�X�rcFdO_pĴ�M��Z��`�Z���D�sQ�_\�JD5�DI*��~����/$eA��V�"X�$���p��ʱ�?EA��Gl��rkC|;�n[��.;�����>4�"۲�މ<G"B(��q70u{y �YH���]��^P�x)Z ���	���e�����y$h�Z�f�Ա�L��?5�v_�������c��|z�&c}萪���\�D�\��Ŀ-�W	P��pފ$M�S����&���n�^��P���� &�e�R�bl�	���:Q�ǵ�݌���(���zt��
�`�zN�#�����o3yϏ�,�u�>-�܉��Ip����q��t�Y*�ףw�<�%�Ɣ5lf��Ak.���Ƽ���'8`Me��T�4�u&�@��O�W'��s�/�����G��D��=f��u�,E_Ʀ`$���r!([3>C\��F�io��I��*���x}��,B#x'*���o�ȗqdg��0�ltWs�)%��K�t�k/�	�o�-3-�Hh�T�8�9��7<̶R�r�����$m�J7��nS�b#���R�����0��������K�QA {�C�w�	=9S��q���Zo�z�$��7��kɈD�x�3[h�;;��/Z7��n����z��Y'!�ޘ�R�Lq�%�g�/AC�uB�ă�80.�ob~�"�h������)��׬�����w�.Gpw�up T"x��ޑ�l�KgPN������%0.T�Q�r��P��?���+\(���:��琉�c��@y�ǒK���|(���!��	ay��=����i�U�	ȗ�y]�V�qh�Q�§vq�[vSc{�e>L�)]c���(m�\�-�I�("u�=N���9#���\�06`��&���f:�q������ ���+*�>w%��FPP����'�j�K�d��{]�/����ǐՃ�aq����0�L���H�B��מ<Z�Z&\���)�9	����Q�G��=�y*�k��U�}KCe.��K�y��#�_�j�S����3 e5����& �.�+aA`jf�S�T�);�Y���k�Iޜ0)�'�^^Ii I,�~��y�o&S���C�k+N�{�&C�E��׻�wa��"�Z��@jx�B>	����V�OM&3:�`�r��ǩ�2��pb��%4,"�k�d�z��}lO���b_�%����g�3�MxFϫ�߉�B]a԰�wl��̸v�)��L]=�c�%���*��,����tiI���hQ�A}0+��7aI�[CьS�s'5���.�Ut4blI n(�w>q�W���"�����KAKHS�4�V�X�7F�D��tF/ѕ�>�H>��ϱ�W�A�q�ˡ�*C�����y�����3�/ާ�#+�8������g���'w�)�&�����s�Q��K��������sš�0�
�[�`3Mw��Ck��mZLP�ǅ+[�U"u��W��mg�����bh�:�L̸L��76�ŒuʁmL�24���9xN�fe*��(�ԙP���_���V���y���g$:��P(��5j3�nNY|F��
�s׳��p��S�Q�׬���aU=�BU~h���m?nG�)�U=c��_]}�[O?'#i�O����}<�Sm��-�G/n4��VLуJF��߿,BO�*\�u5��.v3i"�G'9��o˔��s]4v��sB��$�����dBnEŌ�,�;�m�q���@��S��M���qJ:)��(���A{,1�D� ��扄�����S"�(�nZ{Ԓ�R��@�ͬ;�E|�t���� L�u�t�O�y�4%y���e�{8O"xe��N�$n�: :i��s�,Í��4Q� u2W;��Qׅ�����3*2P�f9��m['�$��FDX��_L06 ���o����k�*�7�\I�S�Ry�,I�I��rr�R&�`�:X�d�E����������C�j�@��
� ���|hR�u<r�?h�E�� ���KV@�CE�ˎS\����RF?��f�����vVSfg�n��d��8I�����������6ae_�m���]���nX���x�9���,����s,+�� �QK�8|��f�	��/��FV=�_�h��XQ�}i9"�8�z�>x,���i^����v�W�ie�ې���MtOh" �\�eWn̬M&sP�D��ɽ`����tF+�l�Rr1內8��W�/9kg*"�<�����A�����jX�Ҡ�b݊`��ohT��x���m`�zX���'��zk��a�ss���1n�݄���>鬄C����"7z)� �����Ks� �l����z�ʠGx�p��I�!+�x 1TVSg�d1��S�;�AD�`t����/^����-~k�@ѡ���������g��2i�)
�nT,�b%Oh�6�,�!�㕂�Řy X��Q��G��u �'͑>��48�C6� ��ny>��kf���hP�)�\ѿŷ���Z��M&�K���}N����zo����7p���IA����#��N�T�>�� ��	Tq���_��]�y�E1\4��X�6s�����[�wA.4��hF�#�n�g��q%�V�hO6Ѵ� \�s��v�UH�)�ш�<�K���z �^M� |��l�8�uH��N(���w�[��q����}JNS���s %}.���{F�ʶ^,����]�>w=�?Љ�U���qNp�PE4��s]^ݓ;��t�	��j������=䍪t����O���y�Y�&��"E2�x���2J�0��KR���3	1Ԁ�Þ[[%$�Y(�$p><)!��Je�m�<�����/�R����*m�J����/�E�>�&�n9W>�l���:��jC�U΃���?ttm�W�s��`�o�i1���4� 1M9!\�����I��Rk�!>����9���Bd���Ȃ�K(i���K�w��a�{�Ʈ�x[[G"�ܸ���N���SF�[_��6�Xu����7�$��(��w���Hw���Az5�#F�30;�R���Iy�����\�ā���dޔ9+{�G����6��B=,�_%"��~�C�E*��u	����:
���gf1ǝ$��l;���k�1�Y]�V����D�T��Sy���ڠSv@ �f��v/�s�zn�Y@ (7�k����z��� �W����:,��Ӽ�pKP`w\�_>�&��J[�Y7����_��JD�nqv��o�$�Eh�B�[�*�p���Э.t�<���0��������E
cTY�x��m�ٞ<����{� e��_f�FO�'��t��A�)����h넮�E>�vĺ���Y�uPu�LQ��\\�ǡ'O)�d�^R^J_Ŝ��S:�u�
���:���~��G��g�wY����̧����c�Z��J�������=@bp��^�!/>��W�1����S����7�fg)��V#�	g��BVI�jE�"ǟH�a��W*��y�����	��G�5Hi7��Th�DpD�ZQ#k�M�#�|�d�6#,OPs�.���2���q��*�~Z�M�<V�}�"��H0s��j����w��?b��r��k\�&�ӌA=�k�`Uƴ�=�W��Y�,i�	�FG��,�?��}�vs6R�.e�� '{̱*t1UR�,֋6��Lـ�_7��d�;�H�Ǖ�u�f���r)�D<� ��	��K�]���n/K~����ݛ�l�A�1>���T�����R����$�]��J�ڿ[P&�w�\�:��1]#�%�\ۛ��>�eԣ��%o�g�N���� ������)dr����t�����`wq�� ��EBج���`��e��-�)��*�hʳ<ބY�ϥ	Onm�Ƙ��⧵7�b3 l�@6Ѫ�����c�z���;	���-@~R8���8�t����V�Z ��P�*��8�DoR̂������`9o�*ό:��c�U���be#u��NM���Q-:�*����iu�%C
:�>d])&F�)?��#Y]@8���i:�#�Qp��3Q=�I���^͚���"���7��-u�Xi߽��|;[���f�᝼'a*?l��w�����5־�E4K�Ⱥ������`���� �5�]������S@4*��K���Ǫ���d �|������0�*
��3l���`f���O���uI�,�F�l��6��%�� \O<e�'��z�R"97~��Մр'�b�Z�f�i����4l�=�����Ϩr���r��Gm'� 4�r{��X<��{�vU����@_� �#��`Κ�2,�#���,�H�b_%e�Y���/��şʦ
ztL��������Rت�gG�� *O��ջ�����W�3+��EU�f9)q����ds�#
��Я[����-�X�-�X�RV��+����x$���;�2�>���eԀ�(RJs]8XE��zlY�Ӄ�LלS1M#�*Ѹ�Gv�'��r�߲,__��W��" ��l�7�RV�a�"K�x��ѱ\�k�7��m�t.a��W�++���2�"�֡��;)���
Rc�&����j�ޛ0[p�݌!�PFȹ�d�7�JGU�BWK�1{T�C|:b�jBV`Q,]�t�Xƚ>S'���M!��Z����;r�]����̒�F[-U
o\%����0�9�^��=�Ģ�Hf�dW����F�d�~0�,�(�&x�:;��@��M�D�O�Cjޡ-rUl���O��ݓA��0�''�'6��>$t�nU�r�ah��L��0x� o(�_����ױ8�q���U5���T�J4yƢ��!L�T�:i��<z΋�c\�1��8��ky�,�X������s� �i�G'D��D�~��3���O:�W����A��-�����Jv���u��Uk�g�HD�r�DJ�aQɦŏql��b������M���?qT	u�2T�K
��_K�Q��������s�鳵�\�J�#Ւ~�k3� |�o��L�6,[ 6�H���|E��Xփ��9�y��=����$r6�7��n�D��2�a�(�l���A����@�|2U��x����K����$��}~/���Z/X/�k8wn�yhD�
o���V��A\�gJc�Km�-nX���=Ij��lj+ǐ���Tl �?K ЌU�qc>� ���'�����u��u"��}|�/����r�	6=I�F ڼ���[���Ad	���5�V���|Υk�fig��r�������:oW����5pS?z��x��
����[��Y�/���V�B�=}�m�@f��'����@��X����h.J�[L�kJ@�~�Ķ�u2��n�fH���`�,W��2��Ā���]Mf�G%0f�g�X��	�<$ܢ�ρ/�X0�Ț���V�+���CӅ~L��_�a�E�<�|���y0�������RF���`�d�6%�< {N᩶Of߇h�rZ��S����oT�
�-�?��F(���n�Qi��< �j��3@H��)#�!2�طl���1��/UM�m��'�l�V��lJ�U��#&{��B7	�+jI���b2��?�m'��:f�W��7�Ԃ�
䶖  �q��cga"���AQ�޵e=G�������j��>�� V��91����158q�<�5r������n��2u#�]��;�³p�N�S�OM�?M�p1)�ױ�|�O�~��Z���֊š��QP:N��ɭn�j��;:�~�� h���"<ī�(@1���i�`�At�ا7�P�#�������-�jc�˖����a��4���_�;���|
(���rr���P�"ق��^�$:{.�?�l_���7i����Ĵ��������(����QN������f�BW��ۀ����m����й�F>��K�N'6�i��s_6� h�^]�+5����\��/��~* �}�f@��ς�,8�(x7��r�|�ՀJ�X(-�I|�^n����+� FE�l���o�Ծh�YQ�p_��F���A���H7š,���f�;7�dg�߭x�}��V���c�x���lm�6"�pu�Q�h"��#��xKh(�k��ď�
`�+�?�D�v����l�ʆ��ƥ���%_�P��'�N��9p�/��Ҡ�;�U϶�u���ԡ]l�U�B/h|�&��c�����<' ���� �O'����b��&�� 61��aBoH��{�Z/�M�p�-�	�nJޓG.A\%�/f�Y6���0�nI?��dV&K�O�D4�G�<������@񌂦Ӿa�M��<ƽ�ꅉ�;�/��?�f1��̨j��^���N��)���vO�x2B���^�ݡIQ:ԉ�Y�Mʩ/�Q3��{ѥK⫠�������Q���2��!ۈQĺL��s�Ü��tP���@^V��+�1�q5p���U"��8��GÈw_}\�	Oe3�B�ť,XB�$�m��^��Ƈ�Sv.�q��L�}���M�,����4�G(� 4/�$��-y��ORK���sDd
0�v|��[v�%�˳1Z�85���I�/Ø��J��-�E��!"�l��?��Zq����&L�+���g���^#�w²�ā 
`�OHu4�x���֍o��R��rK��DHwh��~qZ��s�"�����˲�hd�f�z ),-�����(���`{ڵ�U��]|Px�,�}�Q�0�Qu���?.<]����v/�K� 6>���Wqg�b���M����eH@\�mK��/-D$��6;?%�Wn�4��ɟ
�Ja4��V��~Z��R���������Ŗ����@����j��s.h��<L��K��"�W|��^��#�%VENW߫���l4����n�4�}�A_��P��芑�ny����D��
/p��+I�b�Y  �X�gՅ/,
�^ [�ğ���@Uۺ�S=�D�,}��^�Շ�ʻ���,�6�*�Ք�ʢ(�JJ}�A�F>�A�l�zg�,G��va�Q(0uv�p/���̻��w�iUI4ȸ� �N�|��K{�Q�v�$���Ok)�ĀO��6���ß���_=��g�(
���ʋ�~b^G�`��ղ�C���>)�%K)�r��\��!$0�g��5���z��Nv��ҁf����S$���GĀ�fU�UA(�=u���������E\h�!w}��.�3(G��z5�8QY������/�ř�'�1Vń���i�B"?X@���0P��6]Oa���9�e��XP��*�Z	ߩp����t��8|����l)l[����*�DN�TLEg��0�^���^�f��GP�p-�V�j���2{u��V:�Vg�U��x��Rh��dv�uz�I㴨`/�Ͳ��e�|Fڽȁ���0e9��r���`&6��[��W��74��v^%��H^��i)���u��8D�wuI������d��4g��rE������C���fk�E ����U��9��ª,�c:&��"\�Z�,��]����e���E��?<���KQ}��#��UO4Mל��$l�޳	�,�61~lH�=����~�R�cG��ا�@<q��:)8�xմ�7%)5�^"�r��7�W�G{e6� �~���	{�9B����i�2��+���q���_�*=���ա�I-2s�8�?�w ��U3@va�NM]�W��c<ġ���mGݙ4x�QuV�^=��J�����|�Q��b>۟cú7����U�r�ޯ!�㖠��PBj��,�����!y�_��25\Q�e[m�8{KK��\��7�Zh�l������)�J��^����!<<	�2
.�������~C���4����,]��[�[ONy��t�&��ug�z-���� C�����=��k߇^0��0�Ȇ�:`��N)��uw��&c5�
 �8����07�s���tڭ��V%E��<���1LP}Ҥ`�|E�{���y.4�jd,^+,`U`'�����7�º�-ɯ*[�L�!��f+�j4�K��GB�{s����d��t?;PL��#��/�>��^��^ʞ覰՟�s��Y#_���\��>~�~m˕[��.�P���.t�����$��Qw�K�-�8��'Ic��PP�.1���)�\��������U����՘n2pT��?���.��"]b�z�j:�����y{b V(�!mW�8��H����9�q���O�.[��������B��I�Vb�y��5�j7[TKn�Rl$Z0���'��\��Q�^�KZ{�=��&����iJG8a�{?Bbkm�00۸+>.;I2ۨe>����K*�7�b�����j}��=�j�N�Ս��a� ^_���A���L��#xxO�����w;��(`Ѽ�������ͪ�Ǝ'��ۦ�t37���@�2�bU_W$�r?�صƫ1��*�=�
xܬ�4evR��؃���a0h��j�+0�0]�[1��T�Mk( �R�](��r%��FLM�l�+��:N�"�J6	(�����ȃ�����[�y����^_�Ï������:eҴїT���IP�"rn/`��)��QB�/�o`ަg%��.�W2`7KD�Dণ�ޭ�~-j��@>Q��+���:���[�;5��i�%߯`^��P4ᜊ̀L*~a"�#QLj�����*��M_�5��n���W�
��e��;��s��SIa�!I�MDO�,��)�X_��P3bI�Per{A�tEZ��/��`x�H�ыՔؤ: *F��� �W.�9�}&qO�<g�!���˨���A#>ٰ�6R)�Yi�h��5�)g*��Se�{k��D#pG�V/��
	���}���)R��B�Q�.��nn�A�|5��,O|he���������� �������R�@ٰ��y0�c�N+��9ē���C�W��N1��,md�(��
I�x���2ӝH�}�	@¬ˋO:��}�ࣉ:��0�_�0���Q����E��b\l?��#@L���KT��v��l5�&΂�-��D��ÍH��qy�")Q-y�zƮD��54��}EM������w={kcŲJ�]K������jk]���e�@U��w����� sz�K7i�"]����l'RxYa��[������Y]ǂhN������I�J��
L
6��
zn�h$���ӶS$ a&�Fy�2c�X�^�Y]�A�Z�wg��@�\A�re����d�=>��Fr`� �cHo��b/��䳊1,8��B	aD��]c	x�j ����d:-Q)�5����F���+�ڱ٨W���/�1d�t �UOI�2���N��g��eÌwӇ���d��ySK4G�1� ���9�0�M�]�j�����d>��eF	r�7�A���9��v9�☯�˹�r��b�����	���Χ�
�ؼ����)1�������o^<�m��._��t�@+�Ë�*�ۺ3i�/��]ڰ�W��O쮧~�{�{8Us��V�݊����Yɪ�/�
	 �e���߶\J�r �#�_��;�}�[��P�g��]�(Ϙ����#�ȶ���Uo�y�h�,P���18����<��pͧ �6���<-��*��� (�{M|�m��#�e!	�M�$7���O.�:H�*��>*�/o~���E5�����w�$:�f�8��M9ނ�/:�+�:߰�ސ]`��!�@G5TW�nWS&��F�����ɚA� �x��B�V?l�1Õ��	���$B��,�'`շ������8��]���`$�d%F�ѓ���������]c�����#�g�N�Q ��Uo�5��x�\6�Ba�n��[�9K��{�^�g�DT<,�H��t����n��)|��qM!!���S��&Ѷ��
]kXLoVUS8�:��E�N���r��l���	i$~��)=��#���X�j'��#�ęLO�Aӂ�R,alY��tLC~ְ��H�[�1���)�.��Gc��(��C:wzʼ���ɖNR�%��&>#����n�^��� �c�N�n�"�dם�K�}kZ ��"벗z����\I��)%lŖ��g�<,	�C���vz3���<������mѦڏj�Ѫ�?��3�0����G*qJ�k���$��Zmz�սS��j �B��d�^��>�H�؊-�%����<ht~!Ca���3]3��1/��w�WnE$��g]�H�AqD�����0[�cl,S�O��Br�Y�n1��
�p�<�%`��E���Ʊ�*d4T�8�����w<�g��t��ΨEof�G�e�!X��K���0%��� �&Z=�v�/���ǅ���OG���7ي��0IC��6��71nݐ��~�����EAz�:�:�Y{x �U�&�!��->�`X}���c_ǹ���m*���~���_hB����uQv�
��� x@�8��uxl�Y\L�\��8h샜|9ٜӻ��w�WK����<�|�9��IҹP<pV���>��C�:LF��R֮ꡪ�n�7J'���rm�#]}�i��m����R!�um�Y�j�g߿]c2OfIsw�� ~�c�Bd���*�ɟk�'�߼mA�`�)[�v�
6�U=��wj�\V��R��:�r���)�����1+�+6��+�Yl��ů���9�}ڞ���.���=<�L_A�!3�
��D�6��s�Zdb��ٴBʒ H2���3��L��v���7����w��?��0�hG�@�ĒvC#[D��"�L&�6�!�n��\?E=������-���yDC������G[��Qdc`."�#q�J�.i �6�~�˥zq�Y��9��d�K�ifۘ|��T�����X�m��9�,�I��T?�m��j,8��F��Nq�==��u�:��_(�Oǥ����jq�J[#�����5[3oL�t2�mL.)Q��qoD�z����&D��Ys�&����fױ�[�R��
ܵ���bC�S�����^��!�Zħh�2>�nd��(�����V����0�k(�(y�(fǐE���t���Bh���{�����>7����Y#�� s����3s�?[�2�ԭ�~�QX!w�x���ݿ%�^������}?��bI,���R)p��`,�*��=�/�F��;��(�]Z,���U�3s���@�H��	�U�p��i���Q����~1��B����K�Q�:<9��<������֐����S&��+L��j�}�Dc���� ^�&�qX���ti�nճ��ھsK��)~�䢴����x�JQ�눙vb!����h�x{�;��VI�P�f;�k=K�r�� ~9k8S�����
+Bk�JO�v8���)	-��)3b�d �[�U����KSeJ��1S���D�CRۊ��a�D�S��+Ef�"�'rh�"�s/��F�K1�:�<���S���u�i��u"����7q�*��b��u�GO��B����	VB���j��;�a*b�(%�]A��0���9%(NL���O-��s�Ae�niE� 08t�xi���烖�Ԉ`��Ew��#��N�G���9���J��nU?����﷙�f�����F���^�� ��v��B��WQ+� �lU����d�}D� � +c��`��� [� �6��}e��݃��o�٣uE�A|�Nώ�s ��GK�: �֜�t�Иh
�j�� �pc��N�#_�˲ʌD�u�w�\��_�2rl=d��D	-�|�LK����x��h��m{%��}��u��aI$�i��v��U��	Ɗ]��C{,���4A�f�{�#�HVz��	O$w%Z#�{�R��{�J�p�?=M����z���>E#K�7���Z�lp��'���e��0y����NC.*X�txR%WE�6�ɫ��>�2�ʶ5�:������a��8���/�|F�6�[�|L�����ؾ^��1�j2�4^�/����;��m���=�1v��/C7oX܎4,��L���m�u��{]v0PP�����.52�g��Q�`�r~���]*���j�u�L�H��Y*�A��|̍�$�Q#g�^��1�<���_%�������D��Yj�iX؜e� e\
��φ+������v���h�SB�Z~zI>�E�����L�U�B_����MP[gGQT���)ވv�l�,<���b��D�h��bJ4}P��I��~C��T�����������zmbpt,�80�ϖ�g�и%�B|y8�$g_����o�i�*��GY�lq
4�1�Ae/�
CXDɱkY���M&%����,)���F~���Vp�1����� j�WO�@�:�S�a�AU�������v�I��x��%҄�ZܦI9� ev@L��AU��Ҽ%�����I�9�Շ�K�p$�E�4�k�s��3nd[G:ր��3�T�D.���rS�B�hи���������(�J�VKT�@{rk̺�	�نRq�t)���R�h�}��䎜�S݇b��$3uFmaZ0��eX��oዯc��4�����y����0�z��f>�m@ú��
;��a�,�\.$�����/�d��v;Z�|@)��v�r�:��ӿ����~�+g��M���Z`�͊�z���
�C��y��QX�q�2��UZ|O���&�oW�&"�gܿz��!a.?��$�/@H�_S��Ȯ��6��(R�N��Mh0�%���A��ކ
ߡ%u�cj�R�fZtssI[#��jK'�	;�=���.@�Q�O2�+� /��(9���ȕE�E�{V�3��0,���dѬJY��U��Ч�s��8�	�l=�-��6(сy]s�E������Y�Z�p�bFami����$�$ev�WL�O�+�e*\�Q���Z���<8o�����L�S�;��7�۰<;��&`��+dP��gxŃae�������p4[����+ �Vu��Q��/�&1#⚿�l�2��M/s�Tͮ
ݠ����.#(�ɽ��h�ؓ�����d��_��^��� $x��I��tdO,��[p郜�-�z��d/����T@�P;2�K�r���~9P���t����	���S�G.	s�B5��ԧ�j��_�u���)�v�t�z������5��T{p˧�W�Nn���G��oaJ�V
&��,���h,�5yߧ�Z�Zi�I�J��.]���XY��c���j�A=��7T��a܊�w_�
����9o�t��x_^%�5���!:mO�O�����A�)h����P�5h,�O�"yff���q>R�h*2|%B�5��������G��C\���J!��D $�ρ-�	��cֺ�_@�N�������d�A��5#7�-D��H�奰"T,n��R�S�b��]��!�w�7��FL��Bi��7���h9����}�}>��5Ϊl7� ���3��@?��A��P��#���.�V�T@c� �M�A�K"�76�?�1u�%8�f��mg��k{RǳPH\�@/_/wv�[�2�Ub���'k�h�ʼ�C��W��&�w+,�Z
*d�1~�1L�|oTS�w�ݸ9�F�䖑J>�T~��yl,����g�
�G1�5TB�d���ѹ(���'_d��	�<2��J��la�x�)�l�4�X�$K�����5���WyqE�d��+W\�S���?�xU�bE��hl�ٗn ԘL<>�I]��YSRo�K�&6i���O��~�h_��Go�#����-�B`���╄�$��L_;��є7���d�V!�e�e�_x��l��:�|V�� ��dXᚆ��Sj���e)��=�9 j5e��Xɏ��5���Y��l�R�mՅ3�)�벁���`]�����![�I��5����D6���<�yZ�!�pQ%��_��R��0k]R�!Pg��y��U���5�PeJ��R��^
u��8�9�Zl�4�|3�;̸�� ֦MM�աv3�C �������s��%�}���K�A7���N�G7*�A�'`l�o`��H�k�H#8��Tu�g����J�W���7n�rə^6n�3�[f��- uE܎�C�M� ���$�8#�I����X�B�G�f(�6�G�&��;|�IS0t�p�;DO�T%�'�*�+ƨ�֍���W@�1g܋�jz淆�h���Q��&��7�I,�|��&w5(�u%�ө����Ws�.:r�ߘ�B&f8f�Tk�Z��CcG�ɏr�+��c�Ƒx�U�Gu_z�H?S�ijOZ|�>��ٴ.���]�9v_����p�$k��1`nr�!���ՎW�A&K�*��z��Ղe�1#i��HF8��e(2I�3��V76�֑����$=����[���ΝY}B�9g��1���P=3�c!��{���5���3NΡ^H��k� ���g�,Z�i�����.��]��ViM������؅��=u|e�+d��n���H����
�=������K�	�m�f6W5c��婤�|O'7OT��ڛH<�(xX�:��z�۴Oi���Z?E!U�zO�@����`����7k���ъ��G7-j�{��'�QZ�y��S����G.g�L%�j
�w���dZW$G�.M{�-e D���� ��t+"�p�zPTy�n��mI�����W��x"4�f�1��Օ\�(v�)c�8��;5ܓ�~I�����q�������U[����lځ�y�/���q��+!�y�}�;3���zo��,8���4��O"�5������G���=��/��k��u����M�+�9�6%��X>���ܤoz����.����[?�On�I��qf��{DB��~��Se�'HYƩ(���]��YK��0�w}7?˾IVߓ�����RU'20Y��{ɭ�Z�q�o�r�E/��?tbہ�� �>�uBC��bV~��KPI��!h��<������A;~�`��<�l-ߚ�2��}։T����c����ߓ�X��qč'i�,��
e�Q�V�-԰K1>XW�իA�}�Ns)�9���D4�p��8	[�T�����ƝXI�J�~��}�X5w:��<&�J�cZDc\zbvN`����;]��!�\ l5ZJ�`�����P�ވ+�r��/��{�t�Z���X��y������>��X���ƛ��4|�h$�"e痙�ѝ�de��|�2T�zN�,E���rw]@
`�P���{9�0�d�-�ߧ?73x	����B�7h.��,7HЋkHV�ƽ1�����`XX�T	�O�d����0U�01�1�!�W9��f̈��K�d����^-Km��oph����@80����Aj���U�� ']bh0�#{�)�B��A��������O��I�9���R�c*��� ?E���@�bC�6|g�C;`6�8@S
�zV��
Ir�i_�g� ��?�T����¦���wC�܁!c�q#z|��`I�a�-��o�Z�إ��/�s��y�W�����3�-pLw�1��ҡ.�_l�P6�Oj�t��u�}��AX��!d��C��]��Jc�p�J$�Z)zu�|�~U��	(��j��4�'�J|��-O9P��_�N:Q�1���J��Y�qd-��X������*fv,�Œ�M����3�����بCx8v'�kl���1�Եw�7`�PǞMuq�	C�ˢ��t-��JTzoO^@D�2��_̇�U��nf��x��4��?L�҄w* ��I�(���ou���kf�`��0�W�E_��M���P
�X��uVlVG��Rw����*)�-57����wV�av�V)�R��O\ɯ�Iշr���+��ī��� (��4UԃzD^�t�F:D/_��䡳�m1�c����)��g{�WH��@h�j�XRWE��}�wn�	��kM}�/ީ9LV(����e[�ق�4�Oz��s����j�#$�c
�
��@[������oX�@�\�4☷�7� 1A�WXx���n&��-�xHW�\ ����$���J3�g(&"|�@�.���	�J�Lx]�?�������H�Cn����s ��q6=
 �.��Nq�H4	.P���<+ВZ�����m����zGY7I�D3��v`�PV(������(y���yW����U�5�M_I�,��K���L⎊3ί�2��I!:=� ���b��^��xJ�H�u�N7�:ʣҔ1�CC����rn$�/�b\��7�Y��u��
��o�� ǪS��a9G3���R��찇�F�g8���Dj�pn������Sy�`�&傍��7���LtP�`ݟ��?�ڲ�AA�y0�r�`��<E�bO_�v��Fy%�%�~}7�$" Q���mԵ ������>�n�Y�
c�_������;�}])D%�w�X@%NZ�!;�[��T�}bч@��e���5V7�Q1(�>��l`��}
�d�Ise{�xdj�q*h/��P3i?2 w��qc�m��x�oN��(~�iׅM���9zKn!l覠Q3q��2��!dN�NZ�4R	{���Ӑ}>R�Q��P-�
\_A���W�b�Ou�֧T�=�|�2�HH��L����V Kli���f1tc�8��h&8>�_St�8'u�Q@[�w!4�2��_2�ʛ�G'/�ܩ��<qG�tS��L:V�0���1�Ifs8�@l�K�#i�0�\��KMO����{�F1��qC!��+�Ή�u����f~�U���h �����ډ'FcS.^m@7V���v\��[F�V�$g�2�9W�|�xe�'J������C����Y,[���a�����|I����6�.`�������V��K� �~�����h� ����� 8�� �a)L�s$^��� �<R�a-,!F��\'D��o��
���}��T��x��k�����ԉC$tb��HR�S���Ә�^~�Z7�Q[){�ji=A�A� ʻ���w���3D2�h��O��wZq�>^��t���(S��.��K&��"ψ�/H��Y?�����=�Z�>�vͣ<�_�u�-o�-�n�GRвN;}��%B�n@��ekD>`>��vuy�I�,����f��@���>xJ���V�}�U���lU�bb�x�bBF@R�!n��@�|N�_w�[	.�a��lF��Ԣ���"��7�^[կ� �eD7\���"V�E�tt�D5�y��f���RS�t"�s���`Q�AQ��pYg	��69��DP\�C�D��M�"K�_�<I�Ou���T	��O���H��Ma���ЮL��^tZ���&I.Ƃ�t�)�ɉd���T�&�tr�4X���Aj��<E�7X������"�߼�h�a��)��/;y�����1Q@��d�l8^�p���Q3;ٳ�^"������i�����Q��.I�	��$5��Ew���}�}um)8��@�����}kV�U6�hO���;Ň���˳���r��"�r� ��&ߛ��p����2�-�z�q�n��b���
=�Og_�ƛDA"�������������s��:||�� }�H��O���a���C�7A8� t�m�PJj��2n��b�F ��Mv��=�>���E`6U	���>#\y4ٙ2D�f^�H����`r�e�)�F�En�NMj��ⴴ�l�[�*��$j��to�$|�;�Y�>R"\j���e�a%DW3.R�}��D_�6@Lm;��?(Jtnu����շ�?f�2�"��zXR(H�"=���˔d��$����le[�+���7�S9�n�;6dJ�k���k����:э3��q���[4V���:�w���p��E,rDl(��Y�G.k��BU���'�N����B�"?��2��K�ux0�r��[�A�����|��b��Ŏ��Ė��i(¶|	�-i�o�P(�at�Bu5�j�S���׋;+Q!S�/�vs����뼽��* �[�����Y����~��������:�f#�<��{��ᠪ�U�a�;��j�d3k6�fN�T��D{�������3
��-w���7��-���n���6�����Ǳ��H����$�6g��v��W�!_�����{��G3��GyU��F�2^^�X8!7T]e#��q��uMs}��\�u��"O6҂�jڻ��.h&>��S���a~T�ؕ�#�M��7��1��:SGv��"gqSL/2?)	��V��B��Lx���O�ۓ:�av��,Z�����T����2�����6��$��m֋�CB�97S�ʭ/���eE����xN/����2��� ��
�1-�����߅��(��tmL;����:�ЕC��M�Vt�r�E��vԭ`H2�4��73N��ԽI�z�j`l��r#4\B��4�lm���|׮CX��/$�C���:8�B.	��ec��W����&�3��zq�4QM^�{6U�Onϐ����Cx���8�9�p� �2��|�Q�菐��9pya�X��@������w��*��BT��h���a��Q����,Chߞ������ϐ��x�輊JȄhC>�2�L�6��E)`m��W�jő����E���{V�+��e�B�V���J�oO�i�~�hC<�τ�Ng{����U�[�7HTN�Kb�3>���x�l�
٦��Q���jDӆ`�UQ�*��6H�l}��3�=fds0�5����ʛ�(�x���x��VC4)b<��<��C[�\�dX2_�:���ی�IQ��_������M�ҙ�����;ް�H�H��8�#2)���F��`I�xmK�9Y�Z�o��k=�Vp!]��(Gxx�^�A��ܩ[��R��K6j�!��4= W�_ְ�G-�]}ГJ@�!O����N\K���Ì�/I�3g`"@GB���l�VYM�?S�A���vOޓ��/��� v� W׉[��C��2r�K�g(F
}B�LTe��Uo�YW��܀�A�հ�so����M������b�@"���h~L�M���Wx/�����j�ᄃ��w������K�y�ҹV�1W;Z�ʘ3,h��e��f=����v��	H���
$;�C��K���G�Ϳ}$�z�s���P�t�u�O�`����Y��-a�$m�.?/Y�~� �&�j���|5G� QH��#�q�ۇ���q-��+b\�3�UU���i����$۹ǅ[̸��x��T�ށ��?U��7��a)��J�9�2���Ӛ?A�a�"7����E��䚕�i�U��_�Q����!��6O��>2��%��^�h7�kR�1�5cB�:Ĥ�(f�|��h<BR�hL:+ap�G<X����g�L�·�H�O4a0k��h2��.�dK��+�e�����Y<$p���Zٸ��63���nSU�J��[�2������Zv&�ů�ٱǒ9ΦS�8��d�� ��5���l)�I�"`,�+s_�+��+~�ť����������\�x�y)-�*����g_��ti�wƿ��<h�8d����M4�U�⢼`�&�gX�p8�?!�?���4�&�V��V\N�#��d�S�$���7ӌ�4?F]����h�3��(7^��j���\8���a��i�4�Z�_�Ztq�/x�C��&稃�N���@�"|���a�J��R�]���`�#u1^�D��=@ �$	tѲ͝&?	?*c�2�]�j\�=��oe���(�;,4�z������~,��XK�4��a��&NN�b�������e�e��bI~ �Hw�!F�PX�mS`\d�J��G&�qrr8���0
���T��UwP��t�K���=�:Jrp-Y�㽦�w�b@C ��,'�zC����V�#߫�j��T���l39D����;��oP���{�<*� [ƫ�b7X@�TG�G?e1W�Ƿ;7T_bj�=ۃz��|3���ʐ
����*Uu����ɿ�)W�����oe%*��y4H���~�^h�i;Ƨ��UEd��M�KU�N�6��Hr����x�T���P��^"�lw$��I�68�`%�\�X"2WC��?�T&��2�����y8�c�n��0�>W%���Z�#��"I1�+N
���i�+��'s3�X�	�ҁvmƫv]iOp�T�~-�}�M7s�f0�P����Is��U������+~���I��;�_��v����$*X
��c����� %�0)�zZE�)B�FQ�)���9��#��d�n�p[(���+��B`��N�6�|%3��-G�<�����VA���*7,�g5t��΄P�*?UV��.A�媙ڝq�RRs/��m	Hpѣ�T�zam�,}zu����Q%Y�;�(]�L˦q)@D<����9��Ic��u^j���n���p����R��x�9ۗ�EV�p0� x�]�
���5��On[��-F����
o�x����ᣐ�k��h��
T�%�fWH�m�O��\U�����y��8��@8J"FN�ݖ- �����|�nV.����M$�����[����W���9+?��n�S1�_炵ɂ|<��Ve�q�W��v7�[rKt�x�2�>���q0z����?�
X�O�P�-r񆚹���L{���m�~�0�v�*�<y�Nb���.xq
�FAIQ1���� 	4ЛwI�H��z��VTv9oU��_��=.�W�r@;6a�Ϫ��A<j����ȘY�)���g��)`?�D^m�2�xS������k����u!�j�;�N���3�B8�OQ���8�ͧ���X��M|�j̄��(U,$ �qp+ 4�
��O�%o���l_q"&Se�X<���``̳1	�	��/P8�W$��pL���S��̿�qp.��>*�w��0�m�P�kU����n�9��E����&�Wȃ���X�c�~�T�t�bQw7W�b�Pp�A�ߩID��Q�^	��D�DF�̸�g�.$h��ß:wqyf�UM���j%�f24���E�����׻�e�\��T����r�Y?^]�M�
�e(Xݾ�1�w��X26�������vd�������/Z�������z�����Bj���x4�i�� �"��@����(��s���tq	�4�-���n�d��J���_����ːk�*?N't�����bnm*����'��r����*�]~������k� �q9��Y$������f0��v$� �9�h�, 8��G�G����tD�8����)�����7V�\ S#�'G��v�	�dWL�H���A-܌A6蝋�D���71���e8~��Rﶗ�������[��bD:��]F������BT��>������x���v�N���E��Ҩ/�on���q9��Ce��K�v!:m|���ǆ�.�Z�c���mnД_NKؔR�1\�3\�Ï$���N���}�6Y6�0�`�
�:w����I{?��T�S.F�
:�cv�Q���F��3��$S��Ս�^��~�!#SAQ�3svp��\��Q3^�2���x��rpTǎd�E
�2	_�?mhʈai>�ۜ�AΧ���-ҵ��w˥jn3��������y���&+��LX9��%2r\=�R(^��ر��`�*��l��Gܔ��n,�ܼ'�`�Yx��k�"7��P�fU���)}d���:W���n�H��B%eDCVJV�ܾ{�����8�+���y>d�ɖ�p4�Pg����[�m,�m�H,?$��hu�B���$N�"�~i� `z`�R�$,�(B����^���c9y���H��@G�)"�T�2�Us3)JɺS�͊���n:_�YR����yŦ����h��v'���������KaB�Tw��AJ�Q��X�R�xF��(�U�R������V�ݾM�����l�p�)����Rǆ�ٟLg0��_�
�e�w��6�c#�k3J42g�KˋJ�5~���;�a���GCf�Y˥E1YTk��+�&�6���O?Y4?�q>�.d��J���qq��de�*y��}����?u��3p{l'l��SҺY��1�y���5���	����N�j�M��|�+?8���FK3�&��;���苄���e�9,��@s��i-\���H#�~FxǛ�����ۤ�⦗��󿵕W��c���.~J��u������@�iV�uڒu�/2j�c���+������J-���8)����c�p���u���}d�z��.��Aϫ�jE������+x^Z�(�7���?5/H�2��	���Sr!�^�����v�jY*��q���~�`>������Gz[�魌���(�ٸ��7�la��-�����L�P��+�TI��?��)���I*n(<�N��^F<$j�0p�́�d�b��v-�Ѫ�
��w+׀&M��A���(��s��S���&�p�D^p`%�a{��F5�O�ڵ�:�	���H���� 4������bi$u�Qf���&�S��ԣ��4A��Q��@&�
P�J`��7����j�����R��q����D �3���>��Wd�u~s�_�^E�=:����xĻ3,Q�I+�S��=(-:+�+��j�Q/�HTݲ��2R�7*���ڜ����p��9�b��Nz�}[��9N~ 9�D�fд.�*�ۥ�����K,%��%��id�JD8��ݍ��pB�@�w�B{۫/�.�c�հ������q3���! �Aٮ����x�/� ��C���޸� y����2�1�@��Z��;��r������kED�geSF����C���Ku6��ڻ��H��U��nʯ��8�@ >�1�)���8�r��j���E"��U�}��HX�w��{Sb�������?�dZ�4�з��g��A|f�G�, c��ڹ�l����|]^(��Z	f��>��=E�~�G�WA����y#Փ*g.p���������y�pX�l:#xfs��Lh��Q^oo���M���ܱݤm��f�%jg�WE�(�.DHS��i�yO	g�H!J���z��YM�A�^�_��Ƈ�5�4�j���ø��f$ɩ�*�,[H�����8;����88�()̠�{s�>!+�V���b6keƷ?��S�gӞ�B+�1f��z�}��"�*�V���R�l�s$v|_��6,%&�x��$�5�.��,=�͊_��L�����`�`�����7�T3�"Ձ+S�1�����e�ǥ�,X~[:VMԍ~G�3���K�?�h$���b�:�; 2��J �h!��M]� U�aF�$���F���zK�j8�p�J��5��v@�ݻ�hc7�<T`�o�Ya/&v���4�7Q �������NM�E��/N6���I��N�5���S^���K�`i�j������;"N�\D���W���}��
-���PT� �j�g쿉�l�HS аK��!������֦F!^f�X{d�M��}n�Q�=`tQxih��TT�&$�Uȼ?�t#��.�1�ր��6a�A%�Q�]i���;.M%��S�$6�.�M�j��pܪM1X�_�]�C-ɐL9J#Rd�{���[�n%�{;��o��>��?�&WYo�l�2������w#*���)SUnV�}kFU� XV��f�����lHqS.�vr�b�_T�3�c�6$$jȜ0��2.BR��vP����?��ޙ.�23v�{O��\�7��J]ֆ80k�X�a��^�-|ڿ0��MX�Y�g��JP_)����,+�~�R�ȹ|Z�f� �Ȉ������B���&iM��D��(�Ldۻ\��2tS�X/��7?�`~��A��$�vZ�dz�Y3��#��ɿ
��RĴ&����q��:z�N�v��I�g��ׂ�N�`������������|�i�Ŗ�`�W4�b�e��tu����Һ1�i�x��ȊYk)q�%�%N�'���`�P�"�yD�	�2n#����F�j L��7�?@�$�G��6�D�<���y�֩���i��G�B,8�'!m֠I��Bԉ^H4J$�w�fC	%��N��+Ǟ�l��)��~�fTN����0�e',��1��r��/X��U9�c���h�Dʸ���$fmIY����nM<L�m�9r�q�Z�c�3���Y� r4�C���μ&7Q��	k���r�SCj Dh��ұ׎T��pfF�"#[w�`��^�tP����o����4K��t r&7 ����t�6��q^$֖}d,-�󶚉���^�2�&�k����8爐�.�������W��,]��B�`���/�S`*ߩ�@������4v�����bgk�9�t�`�V��V�������F�KVݠ���J�h�5ƛݏ�xk"�сS��b�ξ�������˝`�K�_�g��(Ҭk.I�j��|�M�!L�������aA�����[$�!{Ħ� L��ҽ$�Ȕt�w��/� O��(��DǼ��g,lc��X��rmrd�4��c�)���ޛ�Q4Z� �_*Ҕf͋䝮��Cm��$'L�$�i�S���S�_RԲ�.ƴu��WȞGI8w�ԣ�9�w5���9?�M"~�w�<���W�8��a��U.�W�+��fZ�~�=���!�d�	4�>OH�h��Ao�`���
}�P��/�v�M���P�In��B�&���˱~Ñ�=���4��1	��l�5-�2�J�7�D��d��ye/(Z».x����yDȧ���V4D]�P�ݫ1����)�����ޅ/}0|���	��ntV4��L����}����G<�8;�\�\$���<�p
��U��8����oѮEg0����4%ݕ3�4�M�Q���$�y�`7,I�
�4(��mژ�S��Ƶ��枡{�*Eَ�Ew#������!k\�A f�&�iWן,�9�Pѧ�K*\|t��NP:�=<q�C��*1}�gA��s�Ur�h��k�Y��1X�E� ���p@0�;�l�7y�u��R֓:z�C�Ҙ�n5�5�,G{��p���P�HuV+��-�1���C@����.�D�l4�~��@/kVSq���-/�p��4zsL�Ox5�,yg�s������N�#���m����I�=<�Vn㖅�e<���&�NHq��������Z+�:��>m5
X -�D����L�3��)	�!��ᢈ�D��P���F���b8X�~�d+�8�>vsXuҐ��,'�-��u@kq�9H߾((�)&W�ܻ�Q5S�T����ڡ.�WI:�v�b���,��:S����M���SD����R�Zqz�!�A���Wx٘4�qĘ�!��qnp�,�E������o�A�ɣ�;:M���H�7~��c:�.�h+��E�7a_�h�����`'KZ+,�Eg�)1��z!D'0P��8��~ѻ$������ 0֖���{�M�sd��ٛY�E�ILp(x(���Zq�|UcYoQ��̊��xF�y�|G%����� �oJ�z����XyaX�����m~L����p�4	|��[]V�*�RX�ޚ���fT�{D�3`��aU�����|�1��Υ1��A�)�Fr]%��������٤���z>΍z�cV�(ڠ���Z�3�#�[#�܏�RZ�����F܂�c;y~D��ܱ߷~�ю�	ď��e5������M�#ޘt%L0^(���ˮC�C�9��rk}Q��[s���)_�Ԭrl�4��E�H�j�\�4���d[Y������@9��1[�"u."����6=Ӱ�u$�P�$f��� �
u}|Vw`|�<�.�P�Ɵ�'�z+�O��(}�@I������wQ�`(�2���3eh�}�G?/�~���0��{��b��5:�
��`�.��-�X���2�R���WU���7�y�lon�'߈��7�D]ӊ)���n>=`2�є���n[����5?�Y�93/Ը^�A�N�����'Y�^r�T1�Nﻉ,5ܰ(tv\��;�?���[��v�JCW��.{��?v�
�ܚWT�F��i�^ix<w�8�+|��4	+�8��K�����rr�,{���� �� ��Q��z�u����<~�)�E�Z�I�3;�@h'A.�js}�<�Q3ԓw2�Z�~�B�����1t�h?ZӤ֗�6�g�l�j�oc3���;�C�X�M�s�i-k�ȠtN�RJ%�b����Q�S�E��Z�v�aQ�u������lo|��x��)�9s���n�Hp��v�M]�Aq� =Ol�����黍����`��zz���,��m��ǒ� �2T8C�����E��T+Mƪ�ѣv�r��솬z��[�R�7�F����byd6�6�M�8���@)�;��-+�Ѷ7%dA������h,��P�iy���s:&W4�V��[wq#fm�@�k�T�����*0��*����&u��͋1��>fl^���jK�ߞ_�	�O0փ	�y
���vo)
�+b:��ˇ샊閚5>���6��=�]�B��-ђg��f��d�ɏ�۽��BU�u`F���������y��<��m��A�+��X+x=�4? �LڧWn:�h�,����=ܸ]�)��&�}3Zq�nU*D.�%G)Yn6�/�LT���:~���~n)p$�OWs�NVW���+$�s�/j�'�ԩe<���~Nq�'��y�\o����m	yq��E!��=;���>"U�b�����tNabѽ�=����C�NM<^�!cf�9����/=ª�WU�J&g��ߝ{NTP���S���,��.�Z����,L�2"��)%���c@��3Έ�[ͽ5���X��^^*j��8�>n��f�@/��$2s+���k`,E�=�P.��p��1��v��f��V���'���r�[wb!#��Te\Kה�eڱ��^\�9�h��a�����V��h�:��_��T��S���}��)�^q��-_yϜQ��xe�"�#���Q25��V2h�8�>�.�@�%Z��&u�s�6���D�*4�%Y���'VI�W �?�/6O��fd�SI8g�{g.��+XR�h�h�5K3�mAU.�a!���3d�>I\�I�ǩjqycO��Ɉ�WHWh%����z9�-a�G�p�����¼�bQ�*.m��#��6�;IZ�A�c�?e(0��"v��Tb�Nq Qw��z�����´����v��?���B~�ç�Y�f��P)�������n[9>��e�A�b(�V/��5C�1_��9t(Kg.Ѹ`��h,�N���0bA����/P�߇���%�=yb�I��3;,�f&�Z�?����fyG��v���^>J\��V�<%/wǟ�*2(^���.6wz�$n%��$�,�c�����+T4)ۢ*����2t�l�!C��ɠ\&�I��Q�z��_{'�x��A��:��6����EbIHQ��1�����"l*���F���</�,��[7�°"B\��-YA;�x���f0��k/��Q�`���(��  �S���5ΛD��hU��D�*����J`�zrF��d�ޟԇx9j�F�<_ݶ���+��sGk*��:S�l��,����x�/�>�*�H�t)Ȫ�8�а�����H����m6��ML��vnau]g�CK���.œPwa�f��
�[
.=�z$O	)�u8�Xk���s#�#k��Դ��)�4��5	O��x�lcc�woF��� "=��Y�l��`���@�z�� �{�6�]3��q$�� $�,����5E��14�ۑ0?�K{�GF�Z1�͵�gܱ8bV��F%���Y�M[������L��c}K1�5��G��^���=����~"Ҵ���M�J
�3��'&�y���!D���I��y�-��;�j�"e�y�t��6��A�����0���Z�����3����Ci`mJ�~���� %H��`eL��B�[�6�X�AA�E�W�F(#tE�l��S$����zi=�*OO������4�����w�wLT�C�0��� e��V�\Q���-tV*~�F85�[�xR���P�O8����MG���a�~�*
\�bO�ho�\i@֟�^���!�j�?�p�	���Z2~_�$��QyyQ�;�Ork̈*���U�f9Yi��H��HZ�?�±N�h����C �1>˂s)�ɋZ�T����|�"�����;��b�#�nC��EE1:��e�<�_�� �GZ�X�x���0ց���J�ܩ3!�+�{1�č�����	_�)�#M���9�fk�>��2-�>��%�hd��G��q��������z�g7Gv�l�I���y���{�T'�{1&�N�8��`�x��Ax�%��W瓚K�S�yCp��:��*I�VO�����ge�a�Z[8�V�r/>�p�sS��z�N���� ��!I�{��+�TB�5�Ĳ�Ws,�_$4X��{o����k!�D���p�'�/K�ʖm��o:�؉/5M�~J$��3�5V�X��gO�m-r��No$�����y�-��pž���K��1~���| 5�6��xI�Y�l�*#�"m���a���[���u�cc�:k��b�A��@��!��bO�d�Θ�n��w	�7�|��k�0<�&ˍ4`h�p��u��h�6��
�Ü9��	,���b�m��nFe�4��XNpBr�_z�$������������D�Ĭ n�P�7����)�̭�9���?�v�hb�A �*4��zt�TI�W��@S",�
Ī5+y`�D�1P�C���^���� �Q�1�X=��It�8�	�0��f���do��:�XZ}�OD����+��~Q�n��1gj���9�.%�q8��,���^v����5�F$D4�A'�1��WLu�2sˍ��R�n{g�e���@�u�m%���t�qq��n��!�	d'ܒͻ�-���j��B�R�K���:T��Q̠�`L�l����{�I2H��JH�1R1�%|e��&�����K��i�M��n���A���e?5Է6A�L���,5cxA,�dqUtE�ޞ��6h�X��E���_���
��V_�D@j3Lb�<�>���8c�ʉ%��~5;x��!���N;����:�#F�'S�\�0jo��-�~��![��{�_�1!<���r+�q��̤��Cx�At%��<�tv�Wo&1R��F��d=̺���B��:� �9��ę�2gU�h݉f��vd�z�jI�1�.�Y�8W��ia����K��It�Ԝ7��y)Y����QJɹ�;3�ѱ-t��a�N$�Z���r���$>@>'�)#�������e��'��t&��Tk�r�?,ci�GwS�F��O_T�Ǐ������y<��ʻ��234��Jg���q��Q����jCrwq.�����5=�̈�).��*�=v���
g?�s�U]���ܗ��O��s�R��H��	���u�����&�d-[o���	����$�o�M֐Y%��7��9k��
�j�ҥ��S�tT*���%a)a]�4�9?#�Hp���b���ڵd �l�,�!S�a��;����R�)a���떓oI�|_H��w�Y��
�U�ư^���S��l�Ws�r���(�V���Œ�_@���h��{��i$ˤK5��fc`���O�`C|X���f^�C��^o���1�1,��?\��9��V�M
P����A�ڒ��HӚ5�LT�ћK��9��纼v�`�Z�>��[�6<����ksd�dazbG ����Ka�+����?�.���Q��w�gG8x�d��Y5�i�X5J�&L�@���x�	�Y͒��+�D�l1�W�x�� ��`�Y��If�b�}�-�-���T۫*�?<��HȒ:�aPCEgA�����'f���|qL��X'��!�Mg:�*�ٛ��V�,�NZ�d?����N,�_���`$L��h��i�o>@"�����*��)�����u���ɉ�#�J	oag��1��!�q���z�i.�.V���-�3|Ӎi��q5A7�#/
a]-|��J�����=)Vd�E�Ê��6����B/��J��J�nF��.`��j���&.qL���D��p�����f�ZKN��C�Ҟ����aEZ7��x�9U'!����Ιv `7zQ�LX;ОR�夳t�W��9�Z�К�y�"�Žq��� P����G陗�Cc,��I��Z���Л6}T`�n�J0m{d��{a'k1m��� gC��5QI-��Y~,�Dƹ�<��%�s�u&���~VyҍщK�ގ�x�}hC����Y&_��4��%F��y-�"䦠u� �����"��%W�L�+hөֹ��+R��»gnvv{��^$ �ؽ�ѕ�C%,ّJ���i�G��<jx�<XeOU��W���	�]O#��:)%?(�!�o���(u����{�y#(����X4�s_��r5?��k֢he�/`��b/���\�(	��Q����&;AO��aHۇ4�[Ɩ�7�ƛ�c��T�*1�n;.8��?�b�U�w������69e\�d���:XRcw� C�)4B4p'���^I�r�ݫR��#��?���'�9k�ắ�ϵ�\g��bѴ��tĶJE.��s���g�U= ��EI@2�+N�W<v�2nO7s��]N:�B�ZP�0�p� 3��R��v(�~�*J��Z�3����%ϼP��Q� e֡�4�<��ם�31�u��NG;���u>�@7�7�#\<8; ����n�#
�Vn���y^GM�8���z3��n�1�6���b �;�&(�T�o������eя_
3� N`�I�y�)��ad������<�9�i�0
��o�(�/N����7K�ZE�#LG0l�d��/�z%��ǐ@�7gH`�肊9�&.L�|]��~%�ntb����;8�h,��G�o�h;�D�!C�%���y��NY<��ԮۈA�gg$<�ٷS]��;P5���v��u�B�vh��}Ⱦ�섟��D�̵h`����ȟ��w�/1�����Eq9�Jx�9�P���~̼7��S�}�1��[�^���}��(:�1���.��P(���tt6���cb�O�%�(����R �5�6g,N���L("F���l�(ҷ�]�_q�ι� W��x�Ε�Z�#�^��-٨�D,�xz�A��<L�ܛQ"��-��&������7���T����o��B�5���C1?�Ƙ�9J#M�Ϟ+��+%J�P�$��d6�[�������ѱJ�7����p�)|���j`&�P�N��ٌV�]��/�e�߳-U�d�i�W븴�21�4�Z�'��#��ip�=&.�Q�?�n���nJ=֠���O�l�z1	n�"�"�+�$l�N:#��{3M��m|]�#�)g��s������i?���8>���/k旱3�z>��BI��ϴE����Q~b�Cds����#V�4.��eX��kn���i�K�}�[!?E-Ɉ�k�D]�s�w�%�8D�e_;鼋.��['�C�3X��5L?�V)���$������T�ܑs$�Ap���x�o��j��}���rx��)��b�[	�!�J�$�gĕ�G� <�ʽO�x�d�<�ʦQ��i1�=eg	�GB���*�Nz˟��7�����U�
�d}�	�y�D%��MQ�ح��� +�ouR�b ݐ��u\YY��ԗ�~%�3��7��,��_�,[c�7H����+��"�(���7}Y�V� �/�ݭfL��.���<w�]>��uc0ċ�uA��͏F,���������":q�Nf^��=r`Br�V�;m���򾙙N8�TM��!>��2:;=ǧ�E[vO�R͉�v�#Û�G�N 4�=���j���� N@�x�{��ކW���D���X����8�}���Y�����B<��@���c�Si�!�DJ؁%���_B�R��S@��DD:l`� Ij��j�5��	޹˜>���;�I�?_���-�]�Г��k[���݆����;|���R�1��:`+�S�-Mx��3l�D^=����+�˺Ÿ ��j�(=��{�I�K #�u����Z���\���'���]��7;)���	������Y�5�,��>��z���Ҋ�J�<��5��D*�[Ýx��jqJ��-	�>E�1����⌵�g@�߰�z��4g`n�Q��z��,S�jNcJ�|�� -�j���:���C�`+z�Ki�i��"��rUً^M�=�۱���o+�j^����qH�Gl�q�|����������g��J�b�5�I��e޵��ޥ�B-X)�Hv�h�׸q7�%� �vb���'��ﾶ���O�����L]�����Z��$��Ҹz��/]�l�\Ɖy.&�3q��A�g����]�t��������&�sl?u��4�=�S��㿹@�2p��؝g��!�o���."�dPĦĝ��$E���	('���W]�)ݗ'������DxWW�0�@�G�]�ް�C�F�H3��.߇���<�����r��(�o��������;�)��>��`Po!ڸn6oܶ06����M�~�j�?
�l�w�	��=��nO�Vٸ%�H��.kI�](�r���(U��;��bU�b�g���Vt�	�� �K~��!�D|=�̌����ɠ��|AW��Àw��$��!ʘYGW{��T*���H�C.�c�K�N3M��1�No[{�x�p�  ������x�N!��D+� PL&6QLT5�۷�N�
|v:vZ�Y��Ǻ��0�u���9����r��L�=��ѧ�R'*��q�vTN~�*D��rJ�}�2��p�MO	k�s��_�	t.<�y��Q�!Cɪ�����n��rO�� R��1��aH�>�WdA��x�k�����_hͣ�񾱥g�=a������9�T�q��l���?]�bx_�v�-�˨��nC=�����dB�Nc�����P�N��`����|�9��Ϻ�b��g�׎=���D&��_:.$E�L��G��PF�l�lR1����wb���T<��/V-��+�1u]z�s����-C]����t0��u&e��끰_�+�ߘ��J��y��jh֗>�"�dm*	�*[^|E�c���PX���%n�B�}�8r�[$�7��c��X�C1��Jnj(�"�x1��v0�ӣ�Fj��|�'iʋ�tm+rd���*�����Э|�+�?�3q�� 3X�� ^!�%E�T���e W��Û�����|l�V���6�,^��A���H�@���ί��AvW���(��<3�8�Ĵg<__�[��1nIή�\�ט����nJ��**_�����a��T��a�A� ���{��Ie7�;hq���i��C�2��y;E��� �t���3cU'�ތ��m����rS��U�����x����$hܞ�M˭:�B�>f
�ܓ��Dç�ȼ"��Ӥ^���wm|��������~�>o��h���cj�t&�fs��Z�~�"[4�d�>�%���*n�n]Y�{�;��`Ȓt�����(�8��p�~��n������Q�a���S9�~�y�&��2|{v
d
'G��J��`�|GJ/h����'�[ QJ�?�}¥@�$�:m��Ŧ_�z��5�-�M+���2�Eg0ܧ�+��}eV��'`g�mhL�:r��λ�S9��4O4rJ��s:����~0�B�͟B�}$5�vUh�0{�`p��Ii���'k��7�jt<(q�����1͏��O�-\ǞV=���Ú�������U?�=�;s��_�Ӯ`�頚���K�#��j�AE'[
����Jb.���>�M�����[FN��#_/�3��6����~C��&g:���XEn�R�f~'9s�~+��`�R�w�M�tH��ŭ���r\U_yTjM�����*�I��ʆ&Z��0�"��"�Q�~�,�)�4��[��m�iT�Z�L���w���8zD`щ�ΌW��.i��\8���� o�B(4��?<&2������s��/�.T��O�+yq����6�xX�Г�@&����<2�ʂ�,�������'����@��;#�BiM�:.��>X+��˖�'|ѕ�`��N%�%�{�D@b����Rc���Q�9�a9���)����hkb�a3��/ת����G�����6���iY'�`��V��s�����V7nDT�On��H�$?�9�����\m�v}g�5o�mq��r�w�w�y{�#�R9䌳f>�B"?�т�/��)�بGm8JL�~B��zj�#$�u�j����=�z��V�a�*���Y�i�������KF�\�xz��:{�dZ���A����`��<� {%,�&�ps�#)d��\�IB�/�&"�Y(�-{���VME��������ƍ=�2-`�V�͵��|}����J����������7�B�QT
��y�(�(���G�6~]�/{�[[0��!bk�k^��+nK�D^"&0��:�V�����S}i����7��4�ӣ5ux�^��`.T8�&L��� E��k�D��2o��W?�Hy8�-+}��r4(am1���n����4]�6E�����F�z�L�X�wxf�`���O�S�@l�di����3����5�#�(�J��@�x����E�Y{I��*s��x�MeV��G;���y7>�*�\��p��C!w
���pK� yOJ������-ҳ�2�R����^��� ��\,L�:@�bA�C]�[g�"V��!�������to5�D��cp��bm� ��in;wŢ��O�O����f�d�� ��+�"�ۦ��B�N��2�/_����O*��x �7��G�ԗ���nI��Ah<~��,�}���J]
9-��R�|�'&�I�}���> �� 7> �N9�����M��Tb[�[���Z"�O�<����H(za���q��N�y�����$Y�����5
c��`q�]J&;���x�MGIL�� ���a5��%�DFs*R�Ͷ���#�l�*@��VsqA�cfL�|U�� ��)ki#��#.H'�/<7B�m;����ק�<�:�%��d�3�_�s�rdxS�K�-��O�i=NI��3�����PncXz��F���YRh���]�i�]��5l��.M�P�����d�2�,h�q�1]���g��������s�1m�61FM�����[��2br�_Hٍ�4���&a����`�M�`qe���ч��T�?l=�-�ݵ��owu�q�7&��ZB��E��t��*�fD�At/-/,O  ��61_�Yc�r�a������0?���s
�Ubc&�#[�#WS/��.�(�%Ȗ���l�^u���Ն�Ĝ��5s��7	s���W��T�G��y7���&�<.WG��C�V������Еj���$	�x�bŭR=%S�hMpR�Jwx��s隔�ȩ]8��ʽ���L�c5:���?�SZ6M�� �M	���>%mk���t��U�����&u�.z�����Q��	v����,YC�{Jm���u���
�٢#����a�.��I����8:��AAv9"��;����*��Tx����#�3p]3�>M�����EP��ټ�NPp��� S�	�+b��#�
%�C	�:7��ƟC�'̄giu%��l>^/s�S���8�#�~��"wQ�DY��鱣����VQ}p��\���I
w��7.�P��.o?�琼@�6����n��ÎE[�_�1�̮	@mN,0s�x���u��to��M)T��F^ J�Vw�@�؎�:�n���{'���)��c�;L�%��a�3��FS7��q�][$���s�>� I���XŮ���`3@a�T��2����1��=4���(��D��������f��KǨ��4�9��6-���\��SΚ���Sl�d��ؼ����,�a�6�m��U���-�p�5H:�ܨx��>�E�Gl�`vq����x�K�3�>�RV�rׁ���T�;�TE���"%0U��h��Pp*|3�����_3�f�g��
�f��sp�)M���1�m���1�fo	����]�����VpO��Zi��r�$�ECh�K�>�9h���Poi�N��q��#;yٽ�W5Qݬ�h��=�&l�2$H�q�HE�YASt�pNu�Jv����3	i�>΢<j�| V �o�����e��Al�ae���d|��꠪:ȏ��sS��QU���t
I��sGB�;�TdYlQ�Q[�n'��k�-bi&��ٙ�.�zlMRmא�e�v��bNMSp�%�k�Ғ�݊��&�}�1m^�|�$0-\�E,��,�2����Pg�$��_n�J�����i�?�u�l�����P,b�%ٲq�7U��M�����;�W{:��a��K�eٍ�|q����c��&!L�X�]�k��0����<Gqm/�z)��@hǋ�x�l�2I�Taxf8JOM��r �6�RH׷�(���n0��\Pf}���(�m"ڑNjGK~'ؚX:vn����5���8�($�O�0]�ȶ����4'l! Mm2�*_�^R�^ˣ����W�����g�5X�:�Q�tS"���=����9\@G�K鮩�:�є�#	��\����|F�s����1$ @��A�	�g��,��En�=td��݊�Y[��î���H�b���9�3v<��e��L���w�W�K��!c�1���z��g��Y��E�\�E���x����l�z�!���%_YuQc��`c��s�@=�+��p@���ڐ�Q_�E�J�7a�	�>���X��P��v[��5�Gsy��a�U���O��7%���O6.+S?�&�3��CwN���1�p�?�
	�B�,9q��xYz���_d:#߿K��������ovq0 i�E�T�}6��a�#a.H�	�0�H)F�vMy����xY�R���c�h��Z~��
z��@j+vG���X)8���A���|(X�3k�Y�����Ҳ�_��_9�.���(��Բ������i�x���;i�@7}�����[7��lWG���v��J�Y�kYc��U���o��4h��Y�a�)���,��������X�i.4�ڲ��a�1r
~�f�y6��3���4�3�3�pc6��۷�¥��}������VE�d^���ւ���t)��y1(�"q������h�J&<a���E.>���r34^,�Y��='~�da٢n0�<��Į_ˁ��!�v+�\@���Nd�]������)`�����	C��0u^��z�Ȋ���{)�ۀ�".(SKz#@� ��%S�����5Ѐt[\�Է�sǂ�V7�#�.r#.�6+��\ m�r���O�̝Bkձ�c}T�u5��|��6�S��ц7_��s��I�Hl���2]Z@%�It�n+|�8�J�,%�ʉc�t{�w�l��aO�9�;l4G�œ{������,g��ƝdEW�oQo;P�3 �}�Nw��q�=��ƣ���4a�&���@��a�؅��Q���0���H^I�|��$�f�u��z2�n�.M��Z*֨��lhM/���acv���<���qa��/��y��Iȏo�&� ��D�ߒ�2�z��,{��L�WO7nE��k\���vH�ϙ��g>T��J���@{��s�ў ��ZBu̅�4C��l� 3��K!��4�j��I�nd ؁L'�ܙ�na�y"ҜI����� ��:Bq��P?�����2�0(��1�U��شvB.�2 Ɣ�}wRM�>ܞ�z�n����������ŕ��*\�sN]'����+͑��|�&�����a���ސA��m�˓LJ	�#�tv�it�V�k�|��Q_"���H���I�w
�u�00�0��l�xU��*�#�tGs��2�d�s�K�5E_}��Λ���~���j �:�2X;m'EM��p����`�)t��_�r,с�(5,D
����1p.cr�|R䑡6etRn�Pq}�(P�90J�A��n�ʓ��������9<���f�+�4XoOL
6�PؕjMj��\�.2�{��\���<2�a�����9��TYoW`EM�mb��1^6�������>U�V�M*Ğ�|��F.��1cfW,C�Ͽ��?�8'�D5��4�t@�	;_�3�r�aem}����t��u�&���3^L�����s_ޚ����hѬ�-A1�卭��rp<�֋&Q�5�%�ް��O����M?�s���*��˅O?f�0��<)�eο������A�06>ƍ�8�J9��2?t��+� �"���0[d�cȫPw�wa�CM��� 3S�����ò�ދ �M�l�v���Y���'MC�:��m��v�D��G����p�W����^�G��J�|six�2�ee/��!�f?�21+�h�K��3����H-�jk�$ӆy����Ri�Q(sH+�/������߁~j�t0?k�!?���us��z��>3��_��OH�`	U��'��<����V8�W�����|���6��y]�@Ӓ�@�6�f���� ��Y�����t�5NA<X^�GB�m�&7)�Fa#@�������`9�*�kwfp�ؒ]w;a�Er]�����Հw����ϢMȞ���ަ��+��s�(H��ܢ��(i[�C
�?q�=�7�LgE�\��.VU4-x�z'�����l�[��>d@A�p��Xq\�l,IM����`%���a�oF���"�J�-�;4蓓�G�a�R���+��x1������Ӹ��L�)?i�	�"�F'���"n�L�������Y����pla����@����2���Jw9�BOP����p�D1<�I��G��)3��lR]�vM�j�~o�&/������){ٌ:d_�C���|"�ڔu\���G��V_e]V�	h	�'��/g���+!=0��/�W����(�xKoFt;��������������l�M�9~���/4С~���Jo�m��n���ny�l��A�<�T���:,���v�>i�lP���x�M/��.j5����D�UT9�(fōb.� ������w��e(u4[>k�^gV�}�-E*���c �U������i�c�̐ �����<��M��c��*Fm���Wc��	����)7�����l3�nh�!�;��+ ���N�)7���T�T��(��LX���r������ܢ*�ByJ	��Â�K6�F��!G�~ӽ� )nw0.�ŏ�8^A�C0��?,���«`8#���u�k��
`�ᦦ���[��V�k�}��k� �$�ǴT�M����Tg��+c��Y7B�"x���BC!���{ �_��M��9k5�͏�P��ѣV}�9e��%��.���E SF_q�e�����2����c��~��J礵�"!�UbTV�Ǆ�����`^ӓ����ޒ�zRg�� �*�t|`��N��d�YfZ�i��=�Љ�$��y�,0���=�@��:�-��;�|�E!�;C'����2�im��ex~&q����Px8�>����
��*"�<���HҘؔ(;���1�B;���o0~����6ǧ��+�c�d������½.r��+�/�\�� {�B<i����JL��z�Yu6*�~�Ό���h�H2��m�'!�5�S�,�8�IG+�Kn�(���+���x�2_-�m2ǒ^>8�h.#�c$���Y<�_,�f���#[���;#
*Km�ɻ>F$U����s8T\����d �=�(Z͈D�0n7I��|l�IǪ�������J@J�� Ds�����
Z�H�F;^���wE%$�%u�a���wɑQ��G�.��tZ<�ۯ��^39��jܙ܂�a��-̉�h�O�>�Q���)�ڇ[]H�n���έ��v��b6�tU$�l����<�~���+x�<���#\{�����|ɘ�<b¦_�U�0�P��ޔ�yCq�;R@�}"*rN�l���
HU��u�c�E�R��?��4�Za�%�2�8&�6y�)qE��w�v��O�8�Q86���_Y)����]?eƳ*q�y�b�k��;���Q)M��2LR.oY���>�@��""e�;DވA�=҃ڴ��	0�	/�KȪ�F�֑a�8�1��	��B�0r�_�'X�c�4�b��׎ݕ`~�`�1U�0�_�v��חgo�_L,㗘$ID�INZ�W.��[�+�e��<B�|2Fy	o���cM(�V����қڸ<�[r��w���t���
!�Q�Ҹ=�ʺ�B����r`�+�b]|da��}�>S�L�j�r�[С�����2O,s:�踋��(�����l�)�7�Г�ل}�&(���#�.)���Ὤ`ן����@xl�=�N��b�Oܲg�ǋ�N����d[i��c ܂�"�c�I���O̫�o\Y(����c}�Q}��JP��?��B�I�����(?�Bpa��X��C�{�v�֕�9q;�yV  ���zC����Yi��I����9M��@�59�x�VǼ8��eS�_"��w4pwM��=<oG������}%0���������`s{e0^`�Lr���NѴ/�$�;�E4��ۺY�C$��Me�)�k�e7�O��b����c"&� �{�'��SS�+$���n/����U�u2u�î�Q����:�\9�2	��e�o0x�A����,R�bL[�<�Ń��'��$�����T�c���B�'n�����P_�
�4����g��w�ꄣc����r�+��&��[��"�� ����e�[�tHrnG�I��<ܘ�;�,%1�Zֲ�&��u����n�F��ɚ�3U���'q�	2�n߼�\�ݞ�8�⡓k#���|�+ڕӄ�R#�Y_�tZ�d�sFJ�\��'-î�h�wC�f5L1�����D����7;	�����ƆzA�������o��˳���JW����R��xB����o�A�+�(89�̘$����k��T�I�~$uc�[��5ƹ�*�I��X�d1��
���篓Ymj�-�C�:��7wv8��v�	��R,�����%4��
�i�2��=�u
'���w�8]bٖM������n������ܸ�n��e4���a��ȴsAw���'KM���c-���f!V���\F�`�D�v�?h����j)�H��Ic+����*+�X�y������
��=n���wd(������N��>5CW��!/b8\=$�F�Xu���zkA�{$��M�KfJ����	�����lV�WЪm�"B񃅢�������Z0�w��o�i�3��
�����g�v(�rw���|	f��' q��qo���^W�<nF�HRu��Έ�զ��۲ �T��A
\)<������-�#�e��b�Mx����g�^E�5�d�3*��	7M]Z�S��t�܍2�Ch��cI�݁K�S�$WF˓Vi���Q���������5E1����7�ɝ9x���J���"�KZ.<�B�?]g('�}���𩡹N�Ǥ����j3K���fOT(cC��xo�=���2�ަ�t�N�G�4���V�?a�V��<���e��5#vg�����a17����X���t��E���J�sAt��c�i`{_��N!L
j�C�����6�`
�V���gaH�V=��/���?�t���4�Ӛ�R���&���,h�����?on��͙�Bh�/�����b��[HoL!_��W9f�ǔ�w�л�j��{�ձQ��3��Vs�����L��1�h��c�ν�{ѷ��.���� lI� g�#Y��f�M�P ^r�wN�t�S����>�Һ//"���!�J��6uEh\�m�/!u=e!qЪ��Oi#�r޻G<�O8G޴z�l���+��Ŝ8 t%��]�v�ˆ����5�������/�����T6�����:�9Y��+�hM��$l���N #k�z���1Tu+�V>ʟ�4D�6�{*��O?F�(���^�y������p.���:���Q�O���\�Ew�8���>^+с�Q��L�����۲&�O�H�����StQ;�cQaԯ:
��fAD�;�XW]3wFV��,���{Կ	P8���Z�R��kÙ7qA�N�-U݈D'����"��vv _��b��1�ÌZ9�c@_��s׽ʞ���+�÷���U���(���X\��*&IX�P�����K�hdAYGY��h��ڒt���T���Y�����ϼ�t|���4Qs/K+��[i�׫��a�'�6[~A��/x�z���G��Ԝ�������9h�A�z�NAk�C���~cy�讣���� f�*�S3N3!�ʁ��?H��,�YnB��̦�!�
�XY猍8�=��������-2:uR���*�3L��O	�J@Z�pK98�)�	R�խ�Z�EwK�]�(*_�opå�|'��m[��S�R���޶��^^�0�8��jd��'@��U?i�!*nW�N�������Xg���柊�\(a��M�x�ei�%(���B)�^PS�Ç�������ǈDl:���^��Up!l��:���î _=�W�V��)�sԯ���λ^8�Yg�/��	���b�@B�*�C�,g�\١�:;�&<���E+��~����p�aP������0�-��y��.��*帨srC�y7��,1SÕ7?.�fwH8U�2��9�ǫ�*�}ܮ��|��]�_�F������<!�>	T���ർ���)N\�eD�jR�a�Szu�}�.��DB�����/m*T�)	_��� �-�{O����&(%�mi�Vy�
n�0t�6Zk�8F�X�����17,�d���x�YǼ+	�5�U��C�x�n�?K�W<��	ֹѼy�l� �_(�F�oDG��k��2�QZ,Ap@�z��$�G��|���}v�W�T���At�I��T6!������@��D�F١��,su�KɲaDN�����x�_0_l�P)�y��P�ݢ��a+O�:/��l&/~���I ��jVw��A%V<$ٍ;Auc&%.y��@Қĝ�V�%K1f��F�H�[��h��8FK���\9�2���r��ϓ���/�_��`j�%��1<��̝evi�$q]֕P]��n���|$v��������H�;~(�ߚгNEW����ebq@�e"9��zl�l�^���X�R�-��|�H܄�!4�3�d��;.*���n�J��SD'�� 2��'|/��"��!m}���lG�����|���Qe����� �����.��0����=�j<�˯��Q��܉�D�L?6W\��Ps�_]̴�k?Cwe��U��<~�L4S�s娦�2������"�C�����<L2�k�M�}�\��/�������0���_�HJ���l۩SP�6|�gvv'�0��I��ɼ	)h�ȣ�Q|Ga�# l���u�G��Qm4py�+��@>|]X݉��Gs�I�r9Lhl�-k��(drK��y��k�_ROac�յ$�E�qL9{����7��������?>�����/�õ����G�,��Á��m�d:�T�k�oТF`W��w����#� �FN����?�I!Ά(�.^<,2NM&,)4�V�>��kI�h.�]�orᆺ��YjG����h^�ܤ�U"�����(tv"��x��w-��@�)o(�G�FɢVK��)'1��^R������=@Ů-��MݍhcFQgv�-��au��V����+��#�C��kJ�x��l���[�ơW��QQ�jխ��!�?0�<#�-�;A�V��1T�(,tS ����s/�<�p}+`6��)���:���2�?�wUDx!2���\;���d>J@��j�ߤ.���9
��U��A͉�؟T�ĔF,�R�_�Ԓ������2���of|z��a��`�D��oi=�X��c[X��3�4C~o
]��5��k@��C�����0��~Z^#�Q�;��˟?>��e`����5�v������z���#�U�E1#�Y��0��@[��6��BB��f7�״��o�R%����`X��|p��W�ǝ�����nt��35>�AËE*R_O;pK������u�ܙ��Ȥ
�I͊(#@���B��'E4���erCL��@�"A��.v��M'$"��x*>�ݭz
�,$K�G,k�҄sp\<�H�pf��Ra�L� �Z^�N±�\8|�״N�L�an��_D��N�
����g>�qE���0���+<rA��_��!m*F���)4��t�gZ�
銻1y�%~��&=3ǙG8�ƙ�Q* ?U�w���]�鎘1���7:�-�h5����~ו ��$�7�:B�0N.}"
�g"�ͦ��{�����O���p��?p���Q�=��G?�_��~Q�a�k�p�MЊ+��PX!�DI�W� ̒��h�L'�����RG$���F��Z�����?%"ʹ��v�e$�����T�^�Ⱦ�Un�'=%)qr�������xE6ӿ�27i{:dܳ萁�zU�|k�{��v��7	7���߮Z*�z�,a]��&�3�����F��nk��גW"���Wl�X��w����m�"iK�t������D����������h�G�����\��'���/ƿ�!��c�)~��/I��<b��q���1�u3��C� <N툀G��aJ���9�,-�V��1�St���k��3�Db���\ ��e��\C���?��nn�8�}��Qo��&�t�w�͢�vP%�Z�崏e�ÁIN<�V	��w�DB�aѓ�Z%L,�Rd6۩3�4ۧ���C�X�ػ)��D� T���'7s��v��l�)���X���ɒ P���z�Q	���኶
�c���nO�T'ɣ����ِ������,��t�
�|/��ʙH�6�t�Z�^��_ ."��������)r��f].x��`"������I=p�R��=O>� �b��P+2�rl���nS��XB���q�֐���� ��ᤇEZ���U����9�	��)��Wcl̜�0��sR���%i��|H�:~�9��7��ZU|�jf����>-6�1
���P����7��4�,R���qwA*�SO��=��[��Y�Mɴ9�TY����6~�ۮ���~ٟ�8;�`!%�,L�}�6��3^a���U_u��Yc;C��c���/@�P�'��^F����ۍf���t5�(�X,��~;7/uP���9�)J5����^�pi3Ī$����Qb���=�p��T^��}sFT}L�3��vQOY���7~Iϖ�Ӛ#�'R���h��c�����&0�芏��Up]I,��MF$2��1��(��l����R�2�9J�V��A�{W�Ӣo������V����jQԄ��'���p�-Gu%�q���,}wy�\�(BH�3q�T�.I>w�:Z7���8k���%����|�3��� �f4��R%,Ŧ�@|�k�� "�_��Ϥǆ������D�<VӐILK �	<L��4���h#��-V��e��X,4����z��+����L]�oiq>{��o$K�n<ʮ4βf���Уi�D�ƫ��o�ZnaѤW%�G��2v�(�2�mz������*��/�o�75�!�Yp�5��P���t=g�Y���u�L�g��k�- ��0o�ǅFu��E�����=x�P���ﲨ�b���8c��b�x�7ӥ�Q�x/�����Ғ��pF�d���+r^P����[:�n����������tr��f�Flㅎ��
�8�Ӄ/�� ؤ�'1 A<��<W�g��6Ʀ|8��W��y|sX���]*�#�ש^�mNѯ�[��z�A�"�2�IC�6ɾC��t��q ]I��"�fm ���~�]c�!�,;kc�2�QW��<W������+��>���
⬔D��OC�~;�?�1��oGK��o�0j��ӔVrآ
O��K��E*�s�)b�%�#�6�YN�ǬR���}��ld���!@Ơ���^H\���hH�1p#���D|\�8�c|� �ݒU.��7\t�}6w�����rw/�U���n�M����s���ZI�����̕�rb��{��fI�Xo!b�ƙ=���a6!&;Cj��?�� ��6��DG�J�uk{�y�_`�*lh������s�^�{�ֺ>�u��)ΡxH^�MÓ���;7|���~�Q���u��uM�%�R�U�~,E����/�0o�P`��ƴ;c���=pL����'��K)��Ԇ;���nu.q��1�{HY6�S���s�lM����mw��{�*h� �i�F�;D�c_q�P�]@���ˌ�>�D�qCMe
q�͙�wDz�U�G�¥���Y_О���`�q�l���R�q*�6@�T�D��S��m���%Q�3x��w0�b� ��A]�P�>�Z��gvm"y��Xvܧ�A�MO����=K�)Q�aT�T��[g�'��+HF߈ؑ ������J̡��r�u�e2|��\{^�L�ŧDo�2"�\��L�ydқ4U&'~�ԗye��؇�Lf����H}����m�a$'�?H��ʐ*X�"i�7t��A<[M�Z{�9�7�Gf��K�nm��@���ӊ�vKA������=�*�CW��|�7���"��-�� (n��m!���%i��t������R�%���ꖦ.].J<��	s��󒇨nHP��܂9E@ǫ���]��U{qT��O�˾��� �ѥ�uPS3�$�H��)-'?w(��"|�EY{lC����G�02�����Rs����Q@1a#����^���|uN
/y|�{�_F G�	HB��.� �b'�����^�!�<� {�WͰ�u!������ ��ٛDo�O�*�*b���ߪ�*J}�洃�m')�K��p� ݂������ ���L�TG��U���Z;�Ëߦ6P��H�z�j1��X�J��0{ѿ�;�������fi�wLx�Q����Vp~�\�\
J�>�?�{|�i�]�F�%�-�r�Z����x�k��d�R0Щ���_R`��&��̰�����ze\�ۋQ�uKǡ�S��Z��9/V���_���QM�f���F�ypK���U
�5�<,PWh�L�g�+�8!�>��gwI�c�15��>c������cR�ʒ�Z��>$%�AtȼS�%��(�6�O�<��{ua�u�6r*����O�"3��/m�<�Wx��UѨ��1��/�(]3vA�n�YSM:ц7��	��ם�>����
��2��,��9����$/���y2>W���68�Hl��7������A��X�'cKߥ�@���$k��_�f=�KV��t6���������_J�n�4L�!��|�Ck/|��L����W��g&��r�,��z��� !���P����e��g�E�)9�.
z@��`������jzV�&���`q��<|��<�@6��1�������܎�G)��ĕ\�#�M>�@�o]`�<w�ڢ��L���O��R��U���O�cW���!qY��y�+�^@��9Y	��!�^f8�\1��Pd���n,�����0�O�1��^�Bʆ_e`gt7�����a��[[ɝ��pd�@�C��pt=K&W�F�t�+(YYα���My�z�6��nhB���>
����ŀ���d�fs�����tD�l��6�qKN؜�~��ؙhe���q���K`��Ё�h���ep��΁s��;����w�v0�i��k��\O7O��e�S�^�Dt��E�	�3��F�Z��rىl����ȩRS����_O�{@w]�ֻl���De4E�Q��ԔMg0�|��U�!�y�K>8K��]OEゴ�A�>6aU���w�I����b�Tߧ`�{%�	4]�Ŵ9f���ˈ��W;'f�TH�5��!l���aK��� zϸ�dǨ
�s͚֓"��x��N��e;Y�2�ֲF8F�P�rK����FhFkB��kH�=D<����^�$��R���yY��WǗ#��Ձ����Ȓ���i��!v��CY*�+��x�r�n<t�ne��w̊x�{�Q���z<k�A"$�*b �s���	;�Z�\߳U�jp�pl�$���>#��?>Ʉz�&�<j3���\���-�H�6�R&A@�Dٿ���'��owj�ݧ;�b�t�W,1lM\L��������9���De(������.�`,��<K��Y^�f��v�%}�!L�����jq�˫�k�Z:��8� ���8n�K�l��f,�ˠn�� j8����(���>/�|��i�F�,��0	0̃V����v�h��CsI�/:���Bn�R{?�Ͽ!�6y�p<7�T�B�g�5|\��^K��v^������D,��5����l�)�>������9G�Iu|5nF/eQ'H}D��V�'���k�4Lm2�	���9ä�����=��Ct
K��[�}��[��a7.�>�Լ~�m���3�-Q���3"R�QŁ�c�+�#��QKI"���l}�}$T�v�+��<�3�4�?!a��O���
�F�n}�C�ʋT��|x���V����m��7�OlG<X�x�w�}k���v�|�������e<XG曉�V��	p`.뻤J�l���;�m�0�sȤ�꿩-�j���A�%��:|)t���|�K����{ ��ҷL}��I�'y�
%w(��tfFbw�}(L�ĔcF}A���b�t.6*f��^�v�E��"�f=�|"�hbČƔ⡖j��x�m��aTE�i�`����"������*��S�kV����9��O f��9�ew`[ů򣜛�c�kv6�`�x ����@�@!*���"4��r�yRś�܈f�l7�+����!8��V �!��c�~�)���M�	�|��6���
ӆ(Bȣ�ܘ�+T�Xu^Mh��j贺X�j}5�햕�����f�T!潨��P `�_&]���$?�N��Xg���t?���q�����(o��W�xsL���<jC,��(�d�O�A3��
���qzu��z���l	�<I1��"��32��J3�T�\?��ԄA�,�U���z�F�ʏ)W@��U@��b�>�ܗ��r�	� @HXR�6M;��l����.tE�"$���(|��dR{�O��,ٖ\$����K�* ���j_|�?!yA���	��ͱ�d�ȅ#�K �]s�v�J������lFS%ÿ�x	}R+T�D�Y.��Av$�؆L�kG\�	��C�|
L��K�ԶX�� ?f��6��	�T��a�9��s�:iQ$��p�^U��������w�db�ѹ���,����M�æ=�ڣZ���-���E4�GB��&?�5��V�ZRQ�;������	j�D���H �#���<y�,��T�����-�AR�\�:�p+�o||��|�D�Fe�}=(�8�����aq�]%��?P6�:<)��U#F�`���~ 	ـ"�r{]`'p�\�@�����3�`�"��BlQX�N'�ob*nAA	F�������=e�ƥ�?&���y���D=�fq�|��X(��[��奧��Q
O7���bXl�oi��:��~J�3ߍ�pF�|�K�)G�Fz�3	��i���{�g��C+Iy��������L%dJҘzC�-�8�6����1�i�P����Y�^2��ɸp��P-��2�� ��:�A�d��c���/�0�'6ęU�`���am- Gk���4�ܺzU��fZ"�A� t����#礔j:̗�(;t馘���#��"L�M�`G4�а�WA൭f�kAw/y�vE
F�t��A�C3�5d]A�Y���&З�$�D"qD���#��;�Ғ�^J{��Ӯ���r�B�p���S�9��ٰ��Oq�o�K���C�Y�C���>X��)�`��XҰ���!V*��f�?y	X,"3�:��X�U =N��vԿА^�;��@i�1 9=���@n8<���w)��?B�!�x�%����������4Χr�j��+O��1[����H���u0�6fq�X�����Eb�Դ5��_�d��� �~���.��>�v��})��d��Q&�{�&Z�.W�D�O��Y@�G��i��)��R×Q� �u昏�c�2�H\�a��ܕ^w�*iZ�n�� �ZAo*Xn�a|lc�J��at�؏���uf?��N�6�5:4w-�Ev7�q�G��G��GLp{H�KQ�:�t���E��H���V�o	>g�@���	<�	���c��RmK����#��������b��9��4��x�b9�4��؄�N���$�F�N<��!�w�=�7��ؿ&Ϯ�#�ހ�裣B�g�4�Tšۭ8��eq��a�瀠���op�,I�O{RJ���ʓ��Bh�_��yأ?�P�+C{K'%Qc-�u�1�p�R�Ғ��>��y��H�\�NC�o�Z�d�@�����U+��r2�#;jM/��2�OI��6~�LY��m�%L��{��Ƅ�ڔZC�T�E{0s�^:�#�Ot�1=��u�.���rIE�������ކ�F��	,���0{Ug�r.Y�F\�?<NE$�h��B޽��X%��+��1⍕�v��p���x�K��@ɭb.��͓�#
� �	���h�B�ށܭ#��(�L��bL�%&�x&i�;(���W6�(�D��3�c����.E)��������7f���~[�A:�`M��e���@��0���R���mq�YG/��G�l �������8TX��ȋ���/��m��e�D�BjH�V9(�����ԕ����.�D���l�T]��>K��1Ȫ�� �n��4&�تi�K�;�y�T����|=T,Ш]�,���R�K� ��*��V���� ��.ʀa�K��T�ؚ@4i;'8l�/����7���Aܠ��4��Lǫ�Ԗ����/���s�����hf��n������@D>\3��J��Ȭ��%����b�8�=���u����W�G�
6�-��=DԮ�A�}�g_�^�b�E����!"都8�=�z�0�y��3Ф��J)��"�pl��Lt�ZO�iP���˧A�����1E��$z5=���#��L>�fka�A"��o��?O��jZ��Gm�eA#|Dm*���囎6��*�h�k�Q��x!�3۾��mq�e�"�U������?���犗�L��F�]!/�5�񡃮�d���r	(;���gB�I���nD�\$���L�����HUP�fXs�I����i�o����!�Y��c��f�|��vk����+�dj~������ɞ�̲*���|oqo�l�^f�j�E����a��6*Wwk#hg��9�~�-�(&�9�� �*>@(q�~�	�/Y9��{rlR��]��DLKÑx��^r���Vl��6gTz^��w20������C;n��Q߳�s'���j���ez/��k�'�?,ي/-��1��P�W0���9��k�a�P�%�S�kz���U���+Oɀo�d�� qp>S��u���p>�;H8K:k&1�j���G��?�����5��.c�����)YU�zۨ�1��7��!��ى[�Ƣ`��$�->��>B��x����& D�|J�Ml�lZ�t��"���Z�[���k���V'�$�*� 胿��Hh�(U�4]P@r�/$�od3��09	���t�5��Qs$\�G9�i�`P?Ù#6�g/��-n�����`�t�
����Ү�]�OiĈg�C��^>E��/~� �vxՑLC.�8��A=/[F+����F%pd�%���T"ߌ8[���n\�&{x&������^�4���Q���R��o2����tu�*F��N��9����,��s&>�dU��zd�(���Wz�����"�>c-��S�2|\��j>X�yN��)2ꮤ�"Cx���L�t��'x�;���	�SD1NO��㔦�Kx��kw��I�L���ĝ�� W���9r�vNdvM%�"\�@�O�Pt=��'�Vk����+$�A�s!�׸׀s8%1����y������	�E@G����C��ɀ*e&�敾�;q�&���ĩ����j�R(,m94��=�;�����%���X�oV /�W�l�%1a�*����h�F�|�F������ڌ`!�J	�0l�Quʸ3������!�h��j�Z�*=��lz ��V�4V��%3&�n��{_c���>`M_�� .AL@
G�TG>�����C�h��fe��br$)T�KT���a�f'v�EۯV؏�iT�Q��������*�8���!&���(Zu���X��B�=��6��[��8�eg��˸����r��	��P�z�3'�b����!�\J����/D��L�ymLF^��w�G��nEG\7�p�m���!z?� �"e��O��Ȭ?�z�YPx�~��M��j|v9V[�n�'�����\�4�����'%o�j�[��R�	�]���yDy9�ᛏE{ɍEǰ�X�s�~<8�� q>Ԥ��u]I|��)@<[�vL��{Ӝ�o,`���E�x,<�3$~6,z�qZb�V��>'K`��������k+�S2F���LI�%
��py�ˁq|eq�6!̣�E��5>�4�5bs����-Q&jZ�HPf1�7�����R���Ъg�P�ٺ��q��"�j�ЮJdEW�_��^��w�����f�����M�����MЈ>�2`A��_�}�?K��S�[��~q>w��\*qv� f�
R�^�_!�5�[�������{Q)�Җ�iV�)�iY#0���K^���}}EK_k�D�b���i�t|c��!ཱུi�+G�P1<�\�D�E���*;hv%~l7�O :��2oOR�_s�r/� �6��O���1e�qAcc�ݒ+TQ9b�0'�*����E�.VK�]�_H/K�EvK�kNk[�PR/w����%dS%�w��0��� ����zO=�`TjԲU����k.��Y��7��d$�~_���h�)is��) �1��A�67��a����*Q���?��Zf��v��cR�%����"��W��ᡏ���DlQ��E�rD��S:H��}Y�U��evbZ�|V)љ|��B1��KP@9r_��`߶��෿޺2wQv���㍉�#���w�nN:�;z�H� al��y�S'F'O!�26��R|��<NN�y+��E��_xڛyg��Fn�:y�A�t��7�����o�Bg���uͺ�u�Gs��˹�҉��5N��6�I�I�u3�ZS��fi�Y̶Z+=Zf�M.5T�,yދӚT	!u�{��i!���d!�;/z����<9X��t±�06"������W[m��:x�o�~�RP�|��R&:4ܞ�G���D<�$�~hTP��&�/:;��e�Q��l�1�Bn��M�0g�ئ7��F��9�#��Ql r�����ٽ��gH� ������#b@L���K�Hl���m��`�!e����5����V!��\���#���\[1��Τ�w$�R2���9O����]���N�I��+��ةg�Mo��M��j���#h���L����JE�Ly��x�M6!�),��~�1������x�5>va5E��d>�p<,����z��zyNZd�?�J	�)����=X�����#8�Vݐ��C��T���;�K/&�qn�P,��5[$e��ǥ���h~×cR���[�O�Ł�n�h�:�R���(¯���4,���,�>t|[~)5��+.ʹ����t�;鷦͊�PI�8��eR�����$c���=��X��Mv<�*��6;�_�Քwpw�m
��GS�/~' <5���Z�P@�1N]"6��2Vs��!��Y�_��F�����s{���!���5��m�N�˵�/�2YloU�>�@����}ڞR1}]�G�%�I�M�ryv��B��ُ��^b)�� �s�hr�n�ve|S��ƞ��&qR�t���_��+c�<E9U�s�?�K�uV-Ou��I�n�Y�%tUr�q#�z�ChK^ܙɋ�A��i��%(����L���"|��O,sU'��_E8��d=�ü�*abN�������g,�A��Q��!��E����zE����L�J�<��f�W'6a���~�9� �=�i5έ��ɠ�J/a�,[ՈA�ɯ��=�\B�j����yxz�P��\kD��Q�@�����
4w���ӥlo� 8mˋw�x���?��m�����%#��s]�uڎc��g+r�F�M�b+4A�|,�{!G9Al
A�M�[Ս+V�p¿�$����Q-���l(+xƘ�f�T8�X���0|�՘�W�J�D�����+J�ϴ�����4�/��(uRw0�>�IZ�%<�[�q���GqQc-���� ��y`y�F�H�'�gGq� �c�mqÏ]���/����}��./���?���\a�!���ԩ�lFx�{�h��y�u�%m!�Y�-�d�U�\" ;��M-&�2�r�!_�n�#e�3��1t[��9���jVn�gI���%��lL�ppÏ�]/H�O�ޖu�e�X�1XB-z�))�fsCS����0
�Ci�D��źw�|إ�|����頳�y�H�񜇙� ��]'�4��ˀ���<����V�.�N�a��kp�JUr0�m;>u� �΋d��K�[���g�B�ԩY
Dh�L��,���D~(�}U�N�ڲ��u%k�o!��⁚�>>B�o����c�=?�ٳG5G�j����TUc�?���ZN#ٶ�)W�,_��.�B��k��r���h��]s�{}�wL���7�}�W}p���4�=l �l 2�xD)��������R��!z~����F�߰�9���Q:35���(YD@��=h!�K~\�>Y��x\UV&������C$+""���(�ݘpu�@k�_HX����|s:6L��7��C˞�9�N�w�]F�Ȭ�U���܁.C��"�
P��2��T\N˩Hm�QM I�X8�%gK��m	�����`�biC������k�ۂ��v7�ܴ���s�� �
�Ý�����Ɯ��&�_iY+fq�S��xv4��.��@�}��
ȣ����~gk�F���(�=�{L	���dψ�i��pI������ǽ��"��74�
����DJ�I"NJ��4��nL:x�|�G?r怃�H��Nu�t��Z&Ǆ�%�݀.|&����\
��ȱ{o�C���m�ԐTU�M�'y�r���X�f4�9*�y��7\Dֻ]��t͢����L���)���z�m���58�+h��ݘHV�ͥC� ��j0��Xp_h��CΔM^��	�=Ӣ��
���k��k}z��R�W\؎�6�L��� }޳�:hp�p�ƣ�D�g��mP��(���a�;�LǶ2���/�g�C���>`-���n�3��B��<cC>O~�.IWR�|��g��V|,P����9q��"���ؗˇ���C��z8�|�?�ݟ���˵��3'�e��*�ƫ������9�z1;:A��Xa��0x��zzw�Mu��%�����P��0P8p��0e3���b;L��g�\:��&pb�N��Y�~
_C��YU9j�]��ϒths���clq�O�3ʎ{�X�X"3�yH�ȝ�Z߮�҉O�J~-t�ZЇ�|������D�̟������ʊ�-M[
��K�{�yy��{�Av�GA��^kPV�M����c��ZD�2A|[8o
�v�,����b�6z�H ��q�G�����.�q{+���0c�?�{75v�
{�������Ȁe����U�0B�y�s��=�oܩ�*Q��|o��Z�t䅬㹴����h!j��OA�3�"�B��*�M�L�ȪGV���Ec__)帧�0���kJ��Q{�(�h�^���s&zAjLA�^=�a���D�9����c�ҙ��]� O�Hq�?��5�&Ѳ��%+Wn���k�W������r$���a�R��@�� ��9�.�Q�p{��s`����uI2U>�	B��z�Զ��mI_��K]46��9�p�&�(AF�2�p��ڨ`\Xm��T"e�a
�O)Wr��w\QCOI3B(�&/&�0i�T�	�����D��I�\\`�~=��K]mU��L�������z+�R�[�$����R%* �!ۛ����>�-_���F���[C�~��"\-�5���E�]�Yt�{�E��ta�ߕhUʚI���k�)�`�߀�x�j�4�h�/c"E��#���A ����{��Ώ�f�;G'�Ҵ=�k�Q�٨���lb��%y�*�46K���aE��$�r�R�%�YH e�#a;�Z���Ͱ�fM#��:����fj����?;^1�rLʖ�n�������vIZ5y��?� �dS��;��žԪ�F�]<P?���"9�����or��Pj�?����AA0r4&'��.�Ѓ�
,-��Z�8�8��(,Ɠ�����^��~�쬓���0!�'�Z#q����O�D|]J,��^���q�<m�]}� ,f��cnB�{˞$�E��ϊ��Չ����p��~�8���ݿ�ߓ�ϝ�R I.y�3o;����%�E��}�C��f-��)*w��tLN<�$CY�C�%A�D���.�w��Hre�q�6m��/����TF.B�P!�̵K�$�_+6���0�~�M�K�����/i�B�N�5���B�g)��܏
I�'?_��u�U�BPe�ȷ�>����P��%���o	������.��;m����>��U_BF���ӊ�[qJk��)X�����Xn�M�J�r��Ǔ�Sev���+�y��>�E�s��{���-<�.FQ_��B�X#��v�r"yIeVP�;�U	�J� �G�g�r\�0�m���:c*�@�����!��5Z!��Ȭ�n��um
�[�kP$�\���(kF�������Y{$�M��}���|A%����5��~l�l���r�<d�פ�n�����:��1����0+_"��
�����[��*���8��96db�?��B7�]�xA�b��҇Mr-�:�tzz��㹽�?��n#��� ��&��5e����ڥm���PT?C�`��`�&[�3�q�*k7�����,U�T��>nPSE���@��>�k�w�\ӿ��o�� �i��I�Ⱥ¹�"Vl���+�����\�$ʺ�m�{L`z�{���>��S׎�u�
�o���t'u�`Z��'=��P�Ǯ�m�w���B��E������s[+��ЅfJ���o(GX~�.\�V�Y#��Xڿ$6�DJ�VG��!נ��d�9O��*�{��`�A�k�E�'�FE>2rd�c0Q��nNA��N,�Aо���zER0. �Z:�:Z!�OWL�sq�go~��?��8t+�J�-�@�A_�����f>����Ӻ�ew������{�"���������g&���㑫� �21������J�[�e�� !"Č�/l."��gN��]}&�&�x�bא2�#$��
��̊�k�b�c��P�FC�%�HM4���?Tj�	((�:�] 	�˻t��qG����)�|�n3����%["dp�u�ߐRH)=#~j�3�J�mI��^Rn�^��L���;}	�a %!��cxA�p�c�%i�g�W�E�,���%x���^�p�l��>�겏�Jj���ԛ�ho�FK8���Fba�Hv�h6�X5�9�C�8 ����z\i�s���=^�?�"ֆ�;�k�{�)J_�Rtd+�JA|��~j��H!j����E��ǌ��QS��D��\@T�3'�7H�"��;T]�\��w��y��󀘲f\ѝc���P֏SߴEe+��iK��n1@� ���*jh�T�W��{�C5p�o���2��`�M	Th�ٖϻ7� ����W���ח���3�1��p�l��ܨ� ���Ԅ8��r����@�A>��d���p�(fR`L���X�O[�T���r���KDA^k�3g=��]{��8qK&�-)
2S�c���+h��=�6{�{23���Y��rq�D�*��Q��9��@��I�R��#�|��Rm�
 ��� ���N��0|�
u�kyf������$�����c6F0Y@�����`L�Q�Uhd���ؤ���p<V>��Z�;�è.��$��<��%C�2/Q���
��ӿGrqkb�ߑ���cL�f\��!��h���D����{c��.Ƀ������'�O��#������WȘ�.,-�	��_��/��Ä7T��!C��G�xS ����B�3:���
Y�����A�]�BsA������4�ZCX5��\�Π� xFf�J_�j�W�ݩ���T�@���!ӭn� �^ M���W�%�V���#!�X�6�#.���o�N`��!*R�o�WO(��������z?R�$��M�
q�Y�@��;�D��4���"��O���%�}�=��m �����\B_��X��U�s�Փ�r�
�?�6FQ ߯�8��O-��H���z|?3(�$�M"��t����R��o��-]}�o���=K-�gEI��
<�|��u�͙;E�KD�)F�G��'!5kXف���hم9Ej�H�ﻝ��M��b���ĉ�6�խh]�������~L�3\/�T�.wƾ� �6�+>$�z���f��`��I9O3E6d2q��Rr��r�/6��R`	c�^d�ݕ��I���c����/��[�|�%a,��Y�G'y�Å t4�t�gTS���9��IX�1`C�`/�U�������JDWH�N�\���v��L��n�/M�O��aˢ<���0�"��T|�WO9yA�0�AƂ���iBck:B� ɀGZ��qC�a����(Á ���7�ƴu[�}�5�����a�Ѵ��p���2Q�)�,*��F�tE�o���U� ���2+������Lvʀ��>���c7���u������(tY���Q��
��͖�.e�^㻑jdmR	�Km���s�U�O�i+Zq@��ҫ���ۉ�7�WR%2 na�5�j$�mW�LT����L�R�1�}xd��5B����N1($v?��~�Z%2�y��y���VCY�7=��`c�f����R]����o��;N��#L��.�/�q0��Ԩ����"��1��2�j�{���6�Ҽ-o������D$_�����S	��C�3�!i�[Fc�����0�(�5>j`�c��e[Z��s�7-Pa:��c�^���2%Z�& b�Wj�N�3uUu"���je;���v�w(sJ�z�aWO��>��O�y>�˨����,*��WU]�1���6��R��@)��Cj���T�����^C1W<_9h����7��p�ā����
��u�d�bi9��T�Lr+�!�ډ��Se#�-r:�Pq-�C��ϋ������RD����>�k� ��2O�Ko˨L��p}��u��7T�����b���oV�(�;6�w�p�(@��hQ���	j���r�����,b.���V_�k�����;9x`xVj��S���h|_���sT��?�r��L�^eµG��)/�#�`��I��c�=��H��re�q�h�+�M���6PSY2�{�ly^>�Ε�ߊ'(�?��ӹ/�i��"~�Ꞌ��\�����\��� �� Ü��?�i��Mj����
]2���E�%<'�Y��X��c�@C`�O��U=�<k*�X��sM��+�;�[�T�h��g��x�ܢW%WLE{	y6��ZIxSb g�i]�����#k��-�xs��kӡ����Y1$��kER�g6��>���?�]���"�_�)���"B@�q"�R�]39j�)���[�p�d�lR\�L��O7p����N4�d�z{8L��͊���+�����܎��Rs���4-�tB�\wiOY�`�|����,�Vo!��S	I5X���]zqHHk��[�٭;��?S��NA!����6�Ϣ�z�	x��g�\�yp�l��?!��L���>mm.�6�}yA�sjy��0ȫ3"�ǵgќ�4f�VR�~L)3�d���Pk���� �t�%|$\��SLL��3��U�l�_�h�/z�R�C3S*�}�v���iQ�E�6���Ao\l��~�yB��Ĵz��7��O��p�9
�9�D�|��Y�!���%�΅�r*�ryƫ6#1���C�K&q���n�$�E%�v_�(�]ZE"�x�XӶ���L��X8SD8����	Y*��I'ϔ*�A YOKK��#w�jh�WC�
�������LLOc�6�QؼD{w����F�����J�Z�V�,ܾ�i�Jy� k��H	K�֢%�ݨ�JF�k���c@���0닾��$�xQvtz��ce��J�k�v�ֿo�&:����e+'���ؤ�55qY{�0~ r���w!�鈑@��?;�u���{��Ҍ���U�v�+e��B�uW�j���ɾ�~����w�s6v�$w�/[t�f�'��Q\�I�dQ���c��`��qV����-8Z:G����jr�cܰ2lK���'�
��ⅹ�F�9���ZZ�A\}Fy��\ĜL��ňH�x�|��� 9���F&�����*Ƥok*���q)u&P�H�{��Vm��'��'.,��p��>P'�oV����#��o����F��@����/1�Zѧ��(m����,,��8�AX���>�iU�/�o��^+9�cX�Mn��� �)9`�Ŀ�}�Ҳ�ef*���C^����+3`�7Q�j�u`˿�����>]��͢�*���)G��%�yZXu��5����M���\?1�xJ�`���@�YLM��5V����x���LR�פ8+)V�RM�oJe��F�@����iJ���lf"�(�
j���.K�Y�8X�J�y5�甡�8�*���O�1�^m)�z,���Y��O�i#�c�~�$�p��
T{ub�(�0�n�&J�� q��	�>v;9޹�ұ.��0;S�W�W۹�����l;ڜ����5>�A^Sڌ�s�S�6��&6�h��(��p�R��Xi�*�Q�ˀ;F��X;U��?F5��O
�|�&?�
C�����H��y�B6G�e�����@�	���-�x}��SrJ����V����|ώuU���	,����2Ľ�	�%í�*/�����U]o�=q��1Fp��)�ܖ,,�	)����T�]��7�0�^�e��0U�qя�������+��Il��ku&:�[S	�ٓ}�J�KRQ���8#�(��9B:/t��,u�*�+��k O�:q����o�(�}q�Z������HeJ�6)N]X���W�rX_��SO`�c�ut��FU(�(@(T�J��c�޸�5�W�� ���1|D��Q�א��
�G$��&�l�����9��!a��!�rN[�E`�b�ģ�ߘ䊍�����o�F4�	�{h�����w�Ř��_a42r����~�1�!/s5�Ŭ3�r*r�c-�N"=|����A��*s��F�^GӠ���C�VAj���AٰH�I�'��mT�n��q�k�����%���\n�w��.��j�s�+����Y��::��/=�dÓ����d#���M;�)պ*�����ߔcw�� �ʲ�h�a�����L�G�P�[�ԥ��;x�}c��ѵ: ����*'J��@��NJ�<�����*���5O�M�����k�X��*c���6UB$@+�J� 
��k�����v�}w;bb�+Kڜ��j��o~�f)rՆ�	����,�b��)�2:�ǵ�
��id89���N�<i(!n��% !�{)m/�o倫���kC���ƇOF�E��b��-$L��Hl�Ӎ=��fb��Q�!u
�����C�տ%��%�O�cKY�W�L����~]���
'O�=[���&0���B^Б�@@��ɥ��3��bUgg@�����Ĭ�8	M���&�Q��ML
��r�*8�ͭTwW`%��D��>3�K
��c�-y�@ύUi[˪%m��3T;Iܦ��5�"G�D��At�	���?���Sd����o��˨q��������R=�6��pug� �N�i��I�����˱�\4�[5:�k)^l����
����\b(Es.�1*J)�ɤ���SPn5E�%��	3sp��Z�QQY��ҭ��b�`��$��(_�M��ϟ6�l��=:���˃-�~X�ר/�l	�hjM�,�'���o�L� ^��1Fզ�K*�sKo2����� 7���]��V��p8>N`�W;�a-e�vw���k{�K�9x�ڄaTt�m�����W׀��hC����4&7 �D�eH�z�(�3�)!�dow*��g�ɥ�r�ºz���[��� i���)�:H���+�"_I�'J�QS)�:�n�!F�;�fM��	O]�\8�71^��A8�A�J8��0�	�"�E$�B��(͆}Y�k�}�=O��#Ɲ4,n����s-}Y�N�/��\1j�H�6��<��kI�r�Ο\�߇��5t�2��*8�7��
@Z71o� \m���نqgD����q]�t�w���9�5$dn/�������;�gW K�V-��H<^��8#�g�u�9&?w�c�Q���Y��|?G��2�m~�c���1���♑�vv�w9�eG��C���{Ɍ>�G�:�4*1?�y#A�4��ǟI�q\��0�7�Q�g�j��T1���u3�
	;P
���X^��w�N�aC)�yE�"�D�I|Hg�`�L;bjg�io
�����J�bo,��I)"JT��s�Ȱ0i?�N���ߚZ��i��������ϲ��3'�V��ٕ�2�B)�3>~��Xٸ�C��������m���1�)Y����h\o-�BK8a�c�9�*Cs��V�U����=c(�z�M���n���~�;�Ⱥ�0Ye���
ϕ`j���T�M��(�y��1���V�-r�~Ї�����T���5�5�� a�:ke�H�a��s@t��\/O�+#Or�(Op�c2��Z����|�o�KZR�;l�A�,:�[�E�~�m5�+.d�_ �r�Kx�=2<)��Κ��\��k�d�z4��zЫ"�$@�r#���Zr�:%�����֝Z�%=�K�t(���2��?3�z7FS5둩���Y*c���Դ��w��/Z��ߊo1�6�q�QJ��-�YdE����L�-�^����c�ĝ�w�4�Gj�R"�u��2'zl��Qq��i�-�L�j(zĞ	 h~�g�5J���+�_/�ESX���}��u!�Kh �����=:����8��!�j�Gp:upg�zڀ�f��Xʽ�L������^�a(V!�ت��"��Q$jf ��PBL1c��KSIn�(d�Ϝ�l��0�+��%�0H0�dȷ��]�p5���e�V���5 �,.gR+��뚼�^��|�l���p�r�v�#�/\�֑�	^����w���eXt��{<Z½Β"\B"��ZʕT��G��L�dTv_F�S&\��Ʒ��/CSٿ�׫�V��1؀�6��j	b*������H߲�Y�Ow���#,z�`��b1+\TZ��1]mo�̉/��OF��d�~�YZ�J���t�q�3w����弻&���,�l]���ڌ�K�����z�36ѓ������`���0k��U\Q�6^0�@�dʍ��^q�|\�3� u�d�x2՝��X��R��TZ������Kb~�i����(�3W���
zN!+��q���M@�U� P5��m�d�K#vT���9[�]4�"�X��{iM*`5[�p+��;@ �O*���urb)�-k��9�^��NnLa'^��g�xWZ]�Lx�_�e$N$���Ma��=;���}{R]Rc�!�ھ ��(�1}�vO2��&�Ok�� �ϝ	��oс}X��#{ǅP�6�&(]F1���dMh�6w��9g�V�z�=Q�J��^�H��}�Ū6x���Y��nj/��<
��M2�DQ2��A���b�7����0���L{�R�q���5�#ϕ���<��8��Qg% @@���$ë�d&Sr,=<w���̢�*w�&���Uz�,J�h�;+�ݪu�Sw� ��R}�o���E�g��a�ͼ⨳����j</(`�%ʭA�I�����J��")�;�7M0�+��~���0�<�B0�8Ψ��#��{���6�_v( ]�KI�Յdn�H�bU@#��i�m׽�ƨ�f�p�ؕ	<Ib,7(^�auVSpV���N^S�/�G����zr��-=����U�#O*�n2�]Q��z9��bc͕M"�s�s/h":}`��C4�z5C��4�,G�u���D�����ō��c�����u(���5��dY�,Ӡ87����ABM�:��6�U�����
`c8���9�ؘ���Ҝ�)���uo�|�`�E�����=I_4��9���>%��h�b�����,K�,p�CI*�1(�zH_p���i2�>|��M̻h�iQab_=}R��	��0
;��[�"}�����0���-[ܑ�~����v�q��w3�0�l���[�(*T6�i�Sm�]R��9�H���B�/%%.u���<��k��1g���n��H�u�Y^�2�*m|�r2������ƅ�� ���$DwHH��JN<)����R�Ñ	 ?f�>�oq0����&�����[ri�0��ӯ�ԯ�2B�I���M^� CH��W�E; �P���Q�f�xpw �aTy���r�΍���t���ff!/STܰ���;S�3�T��kŮ��8Q�j�=�^ժ�R&D�꓍�Χ+�-��Ȓ�xzDL5D�ǎ�m�AFj�2j�]�s�P\�j�����������>o��?-��yB���X���?�<{��1��z@�4N���K&�xf�0���5��p�V�z�d���E�G.OR-m,�9ϱ_�W
��i���N�݋�f��}���,m�l�娻�YJ�ٝ����Jtg�ZůW#)@��D�^��@騭����"�xK���Gm�`r�it~�̠h�
�w�_;�ܗ�Z��޿�����|ʿ���}ڂk۱^��{��˩{���o��Ҳ�>��7hDa+Q�y� �ј�֜�cI_��!�S����w�c]^-pL�x �nPL9,�.gn����^�T�a�?<��T֌눜9lc���>�(ˀ�[V����̶%˚��r�<�i�C����'�6U#Y�
�!qnV�fެ4�a2BB���W���4��k_|'>���D����`��H����e)}ƏPC�����kh�g����Ka'`��TYծTO�A	�~�Qz+aK����v���Tr)֒�P�N�P0Q����t��'�q�?F��u��R%K}��b�*k�҉��y��Q�U����z&mA�Y�\E�� �A�'��H��xfɬ��0t�a tĀKy�kc��c���}I�Oد�a|�=z)�EP�B�GG�xLA��m�� ����H�bE��2�i��I���_����ady��,p	L~���^���u��A���W�Dg��(��kͪ���J�X��xP-o�+����5ұ�4Z��$��Y�Cd����Um-�*7q!����5�ܼ�ԛb/��a&	`�8�6{�� �U�LV5,^���@��@����c�#�h�w�3\#�-����e[��$�PN�vOI��������Ad���a�$IR*�����G�_݄.
\��$Xn ΁όD��)������ca����6r�Л�N��\Q���*��P˪���B�K��@c�,KUf���<�],�d&�m���L{p� �w<_b�Z���m�E��WJ�i��h��=)������CJ9��[��)y'��E_�[}؜z�
69���w��`�R3I�)Rm�R�)�Af��eg�s'�U&)��*��&�0�܋Ƅ�-f5`.���+!����,�I,w����x�#��k��y3�)PNQ�Ay�����S7���~5�DN뭝b(�cH�������C*zx�o�jz�qZx��V����ko��r�1m.�^(���Rm��Eڥ�e��L��rJ���P��?���A� "�9�߿�D^���������r�B��7����{�4�.�A�V���G�9�Ǝg=��(mij��f=�.��+�!o� kgM|���JYSd1����$��L��WU��]�.�����s�1���Ԍ��[���4(!����a^ɺ��U,8j����ON��"td�Ł0}U?��^�޼Ù[=�7���i@G?�����w����PN��pR�QD�),>n�/7tqx�حl�X���z�ekd>U�`����1���]��[ �[�N�L�M9���By�P����O�a�8���X ��OhnCCGOA�2�gr�"��0��#K,�Ef�hx�47��_~�jZ�7�L�^0��^��������IF�D�A�-�j��p~���k�^�m��<���ǰҫ��'�oE����9�gmZQT9�@�U2� V!��~��+c��sB�2��x|ZL7 �ۺ�Ԧ1æ�AD����OV	��v����ы�y�ag��̛�G��9u�Х �����e;������9�ȜÕ]�����ƽj�����.�Q���?ٺ0��1��������#O�������0s�ޠ���(�����#�j'I�)0K�|���#�Ը�M ��N�Fi�!��d��9V��J8j���������4�&	�D�C<1��H�6ni<(�<����9�g�u�9�^A�Hqu�s}� v�i���)�:YL���.(��l!��]z- %�xxV���ϐ �\��ئ�5���:"�����в|p��t�aCϧ17j �@�10��b?�~�n�*�_����,i<���lBJn̅�'0ѧ�PT�^-�?{�vJi��GZw���N���T`��4%�A��?��"W2����Ni<��xSƴ�8}�8K%x�Jc�����UH�i�-�7�3kd���Oc�w�I����cѱ����(sj�G~`��Ծ�,0pq�i���m6o	�Qn;tJ|ܼw�Vs��R�&�2�d�����:X,�X{`��:�Fڲ։�j�I� ���b�`��Y�w�gQ�g�1 P}b��>��L%��:vncR��0ˉ]�:.@��ꀵ0��g��u��y�,�R�nUӗ��$�7�R��	;�=�*����H�R:6i�Ծ�!��Z��(A}Y��r��� 1
�\!� �'Ƥ��5�]�L�j�к#1����s-r��i=�.J��*s�|3��V��l��K=�7����4�����/���ǣڢ2��'1���CsCj$��GW�&n�ԱU9].n���6��֓�AS"��c8��"2����\��ϗ7���v�6D�h�]�W�o.�D�Y��t+t�ԕG~�`�|b�٤���`�B�[��l�g�>Si'�h�4��RQ}��堇�1X�T=ta�|2{r�|Sb[`#��4����O=�!��AOօ����V��z?�������)�egUS��L[���� F__<c�:+8	�oD
c��0�9�`.I-�����0Y�'H���P8�"ö�l5l�x<ɓ�U�:�'��Ӯ!;b�/^T��k̇jm��3Pk��z�Q;F3�YcuA���"�p�O�f
%t�&��$��@ksN���g��F�t���hk�ߐ���W���
@@��� b`�Z�E[��7H�KDFH�)�a�3M��990�]��Ԓ"�?�ՉS�}6g�x�jS��;���c�-^��VV��1�a���3����R�k�V��~GC�:B�{u"?�c�_[��q��J'�_�:� e+˥�=��b�a����ho��b�&�gy� � y�(��\�j�z����K�I���Ç� ��R��|��{�U�r�,�|��Q蜁D���̆0���4ɭ�8 H)��g��vL'��AK��E�d�hX�A1x������ep��e�S��ZW�tI���y��73"Sme�� wڳ_v�ox.Z�o0b�[�Ռ��g��E�e�;�M��8�?򃜰���E.0��A�R��v��j�� 8l'�'[��Rn�ɦ�
�H�@2�� wp_�==��IB��_��Fe[��ʴ��8��ͨd�5c� ���.Y��kD�(��q�<�O���r-�vJqz*��|�B��v)-muO��<'-���1�G��}]��ˌ��I�E/R�x�3��x�������V7�@>���c0�[�2Q!��<�p��T��է��[���v�&���sI��[�
�@N�����=�������;�h��3��@���1iܴ2D)#
K�{�%�ȖND�ҳ�e���
*	)��y��[$ҌG!n�E�(0�GMZ���W{�	�@9��R�2���+n"bjh2F�>������@�`x�������"�+/�4�dV�b���C�����^��gop����A�u�6%t��3�d~z�5�܋v,�M|!5>�L=/�1���x*Dҫ۩��ڐ���lpD����C����M��	.������!�0�P��Ɍ?��ET�0FA�5fn<��	�����XD��ņ���W�5cV팺W�T�������y�������+*K+~��@���Ae�3����gd��&i���*� ]b_���������0������iY*-�����!��蒰�6V@&��ZL�T�:P_��$�������P�̊�C�{��.Ro?m�lڦ����w'�# ��U���д������$<�]��~��+��)��Z)��1�:�X6y�$�zs��L<'�3��3[�5���6r@��L��������a�]��q�O��ҟ�|4��ʼ�h�,��8�o%���X�"���Wbr�8l��<f��2�W���L��:�v�|9h�>�8b)A�P�7���r�N_X�8޺{����h<�I�P���l<��{2 �Oͺ{�/���x�)U���wbwFqB�aw[���΄���Ij|�EE�/}�D�]_j̓��?����:�|���=,�֩�Ǭ��F��H�:��OI@�l^KD���zG�|{�Òs{�y�7R���٠��G��/1 G'�5I���%ފ!䲛.�e�R펬��i44Wկ��Dg:4h�>�"P3�,��%�A����7�1�Εa��!�.�!{�!m!�����Ok��dG'��8��\�0g}�ϲF
���zhΓ���t�l���)]��F8,d_�a#��]����!��b�g�[�.���\ֆ�Fd�
գ��6���	�������:(S+uh���N�Վ����<���iȂF4 �g����7L{���?�`1!��
�?"�Ye�c�f	�,�j� 7�Fy���G�ZCX���s�C��`��\���qo0u��غ���CW6'��¿�
	j�= i`�i:o�J���+0&+s����i��h�=�(/�P<�3Jו��z�J~EZ��'���P�E��2s����7 V��QR�]�6{����l,��,����0썙��'$�Y�Oe�=��C�i)b?�})��<����<�[$�u�_���;q{U���-T���ח�_n��aDz����+\�"��<c�I�Ty���,�jm�V�م�Y�ur]�?gNM�m����a���[Y��U��V��1_�ʽ�.��|d��xg@�>Z��$�/��1�a�*�Ac��N}�b�)��,I�ȝ�y%H��LI��K��LV�-:|�	RR���f+�_�X�#�a�����q9��ځ��+e�˄���ݨ
bK�X
�|�|$��ׇ8u1� 6�^���Ǌv��"/��c�Q��Dc�p�_�rI
h|�Vw��X' D �vn͡�:c����G�{Hߣ���%�b_��
m ����C�6���Q�I���?U\�u���%�� 6Є��P��3���K���b��	�|�uV�)-���R7�9�-*�4�ဩ*��E��[HJ���8����A����y'�Q!&�;l��5���X������|"�1�yav�����n�˧�O����8Ag���*l]>��n\�~���&^`x�P����v��c��d�G>��q|W��|�*� M�m'�>�2F^����Wh〞�Kŭj�W���P�A*�D�=ҥ����$k��<��+��Q;��_^�:A6�٢�뜐3���( i�9]Q����s��%�>1�ɷ�0$��ֹJ�I�n g!4�v�j��t���QX��&&(�`�v��\R�i�(4 �l
���4�'�u�����������]-J�����}�Q�#�#�6D�Q;��ݿA�\�2�G.���Ѹ�'�7$z爘���<ȭ(�$�C���R�%v~�>�!�(7�ji�n����)�ǩ��j�]9�n��H��R�U�U:T^�{�&��4�*X]Q���L{��-�}ԯi��F�� �9������1M��.&�+����0d��.&JԞ����������@�{� �ADJdfA�R�����fʉ�A����ǱYN��X�e�gT{���Q��}�^��|E�U�;~ޒV���ȠT��p5���	�a���^Dv+�%l&��a�}$/\~��J`���,Ti~,"Xy R��Y��@�Zt��c��9�P���5�T_L��� ��Qa%,u�J~K�ٕb�gI��=0�D�{�����́�-�U��@3	M�-ȟ�����{�]h�4���]�Ё�Z!����3���)#	18�\ka��S��@o?�xu�
h%��uiY��Tz��В���b���ԔW�\!Q�F�vB�J�&Z�����
]���PA�юUe��6���1��+�]�ճ�Fw�U��t�˾s):�DX~_�˥�H:wDǚ:38-���o=�
���;:;-�VYzd{�T0y+P�����y̵C_Լ$����Y7��đy���2.h�c�`�*b�%�<�r�qX��S:}�\O&��C}8F��@
�4�B���~l�a+���5�=��.�i��(e��v�I�>��f���BVh�Q��k�J���z�Gw�T|�����L@�6l�҇OјC��ϵI�c�am\��
に+\b����i9��b�ik ���t��=�[@Ț�*����O�Q6����ߒ���0�Ix^��P��m��IF͐/���S�c+�`Ĥ4O�U���2m���䵔m�=�F�,�
�;�l�
^�'ʆ��=�h�X_ �4-m=���Ԇ��ÄήS���.1�*ScM"r�B	�I�v`&�s����*����i��u0�5�jd_�T$^��V"�
��ͳ��3����]���ȥ��Aw�L�#��m�﷿��>�s,�ߨ��mJczu����p�`؎���3Pc"�U�y��QĶE�"���- ���qA9����D`��U)F0+]83�
�9�WAں�b�tg�Mr3����%Qv��]�pໆ^�'�M{��J�z��9H����X�0|F�m�+���uTcm~�B���}@�9�����8��t"�v�?��I\�C��z7'0��m*����&�"���*9�t��R9]t���ξ��m	Z���h�.�����&��F>��W�f��4{e��U�\es @o<m{����4%�!�獗�D��6�Z���}eܮ^����$���[�K l��@���3μW��eZd�u��؍����sl[�)�ZIGi�]~����qꚑxg��e�p4�r�6�Q�� �P��׷�T9�Bګ���2h�RVq�?'F�=��0'��D�~��m�������S�	���El|&jS��^��c�%��P�(���~z}����2[t���	㕣wU��RJ?�b�>�:�<s����1�+��;�J�� ��}�9�����]�GE4�hM�/*ō����qMd��ԣ�p���uR�C#�;�O��l�-�-�R�S�����{�"�� �9�^�=�f琼j
��	-�5"\H�]�E�������+m��Afm]0���ήۖ+!�^�>�Y��u���Ԩ�UF��bݙ�ڗ�ڽ�gH�'��.�� �i'c����jh�TU��YD��zF�H�	�Du�Uy��02H�a֡;��/��F�P��h{ȑݮ��=u�-�[����M�T��(5�1pWc��R�"M�e��C�T�f1�l�;��r������螄�Z:��iC@���}�9:&���zMl��ߋ��Î3�M��$��˰N��R龺PBRL��uW�`S�I�1�Fh'�ŗ��Q��<['���vA�;ԌӼ�1[j��L��Hu6]�\Y�a��r�d��N����>�����9漑�5�9\gH��4���Ԗ%6ζ�0M:��Kv'�W^�v����B��\Ya��Q��q��� h�u��i*i�X�9M���d���~�I�Jݷ�e�{���}�%V
��:�@��:L��X���gF����q*�6�X�v#�+K���a+*��ו�UT�I��e�_{v�X�[�}��)�e��UUt���N�t�����]a�	��3"�p���+��� }����7�r�'�x�/.0����aO�&��1xl�#6˱�Y�#t���QB شEϥ-��"�3']�iV����w��sp�G�����;�S��)��ق��ES�R�����aO�B0��Ւn�r�~>p�!3��-�eK����7��J�i��;��%�mc�Ry�	R��\�ʐr��=�!�/�w?�8�U)t�+�H+^�<Hݵq܁�Z �����	jf^Sr�xT@�A�>p=�+���Ff��T?���o$����p;����IɊ���Ah���I1Z/ +k�fA��@�iY��I-��n%|�2"�J	����f���o׋J^�h,�^aIy�]¾��W��o���舡�ނ�R��wb·nƎ������ؽ�|�_'0>��,W�
Z�a[GIő�VL3B��uR�,�Kd-"�tà����=���<4�;��#s����$d%so�V�F�f�M�
�yષX���u�r)-�g֮%Ǣ+��2�@����@�iQ��K�Yp!���࠻�oι�����w��: BW�p��>����q�������,�S�9���������)�>��4��1I���▓�v�m���z�؎;��T_|az�rA��W�{%U]K��J�]�,ֻ�6�/j_��ώ��W눾jE�ו�������K���%t�iH���Db��2��C��!�-��P"�T�4����l\̚.tm���N�
*Uո�w�QP����r�|�^;Q��{��/	ߑ'�Ť��ꑤnI(y�F�W����;�NM�~�:��r7��miz��s��k�Y*y����)�Kg��z��JL�����#
�ߢ�����P���)�|a-�c���*��Q'�2`='�mARۏ�w�2n�ns�7��|�������p����T�y�8<Ĳ�×;~Y#�L2���Ͷ|��eR,	q���` -�w2
\�#�hL�7�*����w�6Eܲ�m�� ���	����ʈC*�[�ngƯ�ַ��ܭ��ԫ�OmH��T���L��"�K�Iq��#CdfZ�S"�|2��R��︍�@/���M��d����V�c�(<]����Y�H�8}Ko�����.ÏO3�_cl�u�:��Ȝ�/,j V5���TT��N�)�$6�5C_����JF3��p�
q�H2_6`qAm�Ul�!x�����o�_�4D�����B��_��J��P	���,���Z�.a
�v��z�#}1�	*�<s��K�0��g�Pv�OV~L�B�Xe4W��PlØ!�1�P���c���Ȱ���31yO���~ w;�rt
�-� �m]�e�+H[��y�,�"d�O#9�\_�(�}�����6�?0zr�F���8�y�)ѦN�k�Q�7�ɪ��.ֹ�z����0V/X��"�QaO��O�ը��7L���/��/ma��G�h�cR��4҂��h2��k��;�R3��nx�|���aJ�X��O������S�^라H�ּ'$�W3^���NX��xng���[3O�hLw��41UOё�ċ��Q�����A>�����\�4x������|4�QDƉ�@�*3f{����)*&X~�nS��
e�&���x)͕��x��J�C\A!2)D���R��?Tv
~}O���Y�e�q�{���ĸX��Kz��ɢ�"c�e�iܩ�Kl�PЩΟZ�$����K���Jx7�砖%[��tp%�pG�S8�ӷ���]��h��~'ƪ��7j�j�D�ټ���(P{�6I]���$���ސ��A��f��9�)a�1屇�,E�Oǜ�Q�8��*F���Oсeu2�r�si���fe�%�x^������X��NH�]^>���V���٨����/��[����7/=���R���\&?�w#��7� �bK<�qϷ[��d�Z+ve�s�gY�kr�d��`�I�N�;B�;f�fS��HL��e�~;�������o#x�7��F-��.n�&��;�]@����r�-���-�^+��?�jxྏ�K�q���*��Z@@�8��R�(��B���/��|&TuƼ`�,�wÒy���y�출�!��F��|��+p��G�i~
��i!Ц3y���!MjW��Hl������O���C���r1�EQ�Nq"_{{��!�����(��+`�J�=#�*�Y�8>�I��P\�}W��Yz ��P����><d'�G�qϓg0'���T"��n�i�ejG�zd�2W�,3?���>�kw(�N4�31���|jS�$A�-���U�h|�Cz([ƪR�߇��6/��ZR���U��z
o�=Ͼp�'G��=m�.�>1P�M&��c`���p��t��l@m~\�x��C����$sڒ�2���U4sIbz&�b�W�7�T���2���dH�x�ƒj8��F�Ǉ\Ɉ���K<�i������*4�ZȒ����8)���<�}����$˿}�����ހ�2O|��Ô�2�(I����L��@��N���_Pp���".�C����D���7=RQQ����ҁ=�6]dS���
�{6e^_���i�h�D9-�\����oCc���p����+�y��{j�#Ӝ�D�BPg"�&L.
��`W�vo\��������S�[�_UswN��f}�!B?H9���x3;�#�턜���'��`]�q�VC�2釿�Ec��38��g��d7:�sh�X������.�Ä:�B[�<���� 3=��O%�D�󝄦�)�]̩P���46{;�������yjJ#Y�ɬ��;X<y��o�:�K}P#���B�m�
��0�="2m��JV�y�YO@2�8�>	��{��t�nH���5h��_�­���.VX��<������M�lq ���V��`z���롸ޭe�Jx��e���?�ޑ��_.� fF��K:&�N+8�R�H�;:�� D��6�ª��HQGRC�(?�ȑ���#�+�y���:=�}��w}�xw�:�}H����	?I@��$x ��v��������uH��U;�c�R��/�?�E��Y���w��ȼ;9}�sLRj�� m�����yhI�.�׮�To60h�H˼��`��T^}�=��L��)K*�Y����۬w��]b��>dI\��t���Ma���<ZVEV7�صƍ��E���0Q�b�e��5���p3��%>��
+��8w��5t�	s��5&�:ng��Mc�N�|�zN��HC?�
 [5F��5m��c�mA���"��Hw�	伽1���ƉrT*{޶9��Vu��q��O�^�EL�n��nE�bA�@gX곜H��I��&�/D��-0�n�\����A��J���(C+$C7+�Q�|��ǒ),�D'`��/|�?��]��\�h�����-�U.r�(�d�1`
�n�4�{�$�R9�k�Wg��03݊�W�	���۷.��-g����i��{d
��H���%�J?�X���D�]3�	}�5��i�=\���v�Q�0~�x���%����Ŋ�y0]`��a�: ��;@3��&:������[�_l[�:��f1	G�tJ�Zb��<&s�r�.仂��ZXp5G���l��4˓,��1袼?�9�^6j�u~�0R��I��T"}A�s����#��[�L���p&&g�\;������A�g3��n���"I�0����9�G��z�}+ǐ������|w���;�$��=<{�����|n�)��Ώ0Q��p"��KH��|4�:)��,� ��k'�����������G�~!�'ɏ͛&�Y�	�]׍ ����D��>!��Fw�ո�R�"�t|L�Ո�wkfʝW�#�n?��]8�:q���qyy4�^��y��d���lÏH��?�_]�?9�c}4���Ⱦ, ��vqڠ )�´1��/-�d��{�9S(`��9�H��r�ZRN�4�>�7/�޹x*����u$���M��_{���֬(ٜ�p���ڹ1�v;t��$��?��������
M\�4���0qBtư���g���#z�z�w��k��V�9�^o����q!���*�11�4�J�̹��dPA7�ea�JdZSm�jp���Fl��	�X�L�6���o?Ÿ�<�vC]�Ճ�,���q�Zݙ�̂�~:�2�Q5�ل�<���w������t��4*�uJ�/���X��7��Ĭ�<�KW��O�H^o��ŷ�m�:�-N�-R��slw02���ֺ�f����
_̠Z	���D��gưV���1Ny�w �c~�d��y����8`"U�[Ķ�$�L��p�z�[x� ���2M����6�EzR��y�t&����C���sn����뗃p��g�w�F�t�#{6S��zO��Xt���G���9��⨐'��������9���\�:��Y�/�7�$A�-?8�n�h��>�'�ۨ���Â%���D!��k�~���
��
u��N����%�!X���y<uh����yH.�zm3}늚8�j���\�lt�F��1���-��z:��L�����jug9�y��
�ALr/�-P�:�C�d�R(�~��\�������IvX���W�Zf��^�@�\r��Ԕq?3�����T}�`���O�wG��	�#�����	�+'����_ou�R�sn�჻���<�a芦��>EW�E8��C=�q�b�D��s\�g�i]|]ރ�N�"zF���F����F������W(�ή�)��	���X���u�]K��Uˉ�4ZBW�֖���u����w?ȯ�/�����7&|�d}o����%siU���gj�!�g9O�|�E[tM�<֤�%��O.6��3{���А���+䡢��c��}��P��
����
�����tkh�k�m�u�F{���g��IC��u�'�x�����RE���~��f�#S��.5
��K��^�+= ���b�� }z�#�t�b5ɑ�:����9rG���W��̿������}�<i-��L�;r�aj��xTY�+�g]� 
(E�a
z��1�q�����2C��i��%!��@�4�2K���V�fo�i�PN�VR�����H�]r3�R�6x�}$��4V���
S
�x��Ó���L�� ��̷��T�$]01����t/�A��W"��Jh�E0�q�����y�,�O�S�н�^JN�\�����@p��݌c=�}�	��y���u��Y���Z�ΆjӀ����d�����3�\��� 5�����Ju!�{�z��V������_R~��y!u-���E�[m �F_/a�D�*0®I�e�\���pir|q�ѹ�/*�A�w�Mq5�+}���B�Ώ�D��n%8p��/��5N�]xr�qE�|��������L�5lf!G�i�}z���V)��0�/��u���-�䟷�M�|C�:"��y���-�����:��ZIqM��;DF��D��gRR�� x��]���.��?�:w#,�
@��׆�j^�2�3֫�`�ή�9��#7-fj�x����R�E���wq�I��\��)Ja���/*i��3��,#T>J0�V��h��nzԫ�5�FA�b�`e�r�38e��/wm�� �:��Z*r� ��$���O�������_�Dv���K3���BS��QH���W�|N�P���`�yϯ��"��yM��)w<�;7��l�_e,�u���Z�J7�43;�	]��+��F,,�T;�-��u��Z[��Ӕk0�Si�I2q3�.KN�v��%�Dlu}��|���}��Ӈ�Y6)=��T/�����6w{��W2 d3���-t�UJ�F�l���I����WUĹ�d����o��Ӂ�	��6�h��+k���^�T�����y�8� ��Yȓ�X?*�6����?���Ȫ�>�L�L�S��8��� Ab��
f)�9hL.ً}��;�ys �������g������:^;>1�b�$�0CE~��/�ڠ�=u�J��Nq�逞�3ƀV3U�͚d#�i450Ǧőȑb�S͚��[J/�)z_ެM�J�tb8NTl�UK���[s�$�QL��²ǌ?U�Ć9Y�Έi.*��^&|
�x�-�}~��?�JW�Qё�gށ˪gW�W�@P��E5u�J�w�r��&�����	O;z��Q����F�x�0�t��]	��H�{��=�������a/�f銫5� ?�,��6�R�ㄇ��Ņ��\�1�࿙��f��K�Sa��m�=�z��� �f�h���{&��C0�VɁM�H$�t�´t����6�e�d��k�܊�錵�o���f	m=��z��a -����Kܟ�AS��LKf�g��W��lD��S�a�̪h��+�պ�! e;��{�D�^�c�3�u�)1����(p�dp�L4��n:
u�aL�G�%��B b1ٞ�V�?kKY��w�]��g������k������~��8��'��F��M ��\�[��Aguc�"�Y��e�Mfl���:ޒ/ѻ�8,���Y�%��Ly�j�,&'��j����l_�EJ[v�(|��T?i�ݤoFޚE9����=B2Y�� +�U���s�Lu���#�}]��.��Z�^I����1�����)6��*��E��EƐ9�����_��0���E#~}�6�8q]�r2�u��%����(�u��ɕ;X����lfmȓgJs/�J+$��c��y)t��1�TF=�[+��IϾ��ͭ�~�Tz�
�{|��_������6�H}W8�u0o�N!�4#=t����+����_���Mb��7H��#0��W���5�{��s�θ3S�fp~ۥ8*�����
��,"����ödJ:qLDO���"4��_��3�]`����VJxb{Xğ�t�/�ڹ�FG��~!�nl�W��uT����N/jmBc��k"��Z��|Cl6�?N_�L��s��R�W0ﺣ�5�a�|��M�sJ>R&A����4c!��r꫎�!�ZTz��_v�ؖd���K��9����A��Ʃz+Mz|�0�0�uW��h��]l��~��g�B~K1�v�?��Kg3�{ge�dM��Ъ�GFr\�V��n���2�9���O��V�o� 1�!�o��D{��lǳӇ�j�e&��J�]౾�&���(��E9�j����d���]q������/�?Se�S���ǚ�N!r9d�M����.���c�Y�,���v\&��g+�cS�c��k� �1�9v�)�i[�x��Q� �@�X��-ϴ��(�V��Le!�Z�fD���RTPDwЩvaa0F���͗(�s�� �p�	�t��H�@����4�nw"����g�$��y֘h"�g��R��^�W�7t<�O�]��Yw�k��(��P(��y�ऐ�W�m�#���6���(;���X�����m,t���2���޺ ���%�
��&��㮹(�M��J�/b�� ڦك���}�Km��2+C_��?��yt躖������2��N�o��2m�J�*�{�^,�p : ���Dg����κ|\r
�-i���)O�6&c�;��u����'��0�@��x�Ƅ8�:� .rR���G��A֓!�0,.�m���F��{aܡ��jL�jس�,vw%hE�p�����$B�8��֒7	?��==�z ~���Кɹ���+r��1��w��$�c �Ӽ���"jt�a��a�ٙ,�����AJ�Ƨ�dB��H����6���X2�rQM��U���3^����{^��g/h�,ROGo��h>uod��v
�I�]�Q�sys���h�1��a��	��G�RB?EѧJ׿<~a��GI��NP�����{�D]� ��hJo�����k��F��ANW�~5�,�O\OH��
;T%U������!+d��d;�1��X J�~�z�/�o>a�U:3>�4u^MP�<S#`�o�K32y+��;o��
.��%UQ��<_E�k����?���6t�`\� ���nk�d �:I��}�2�4�?i�x��f(0����O�F�fH�t�G��{H�s$+)^��F�����
�8S0�Q�/~���r�B�BɬF��d	�)⹩Ɵ�EVίPή&��}>ȡ/�]5
٭?��#���C���/W�#M� h��g*��Z�mԎ�	�"P���|>2 �K0���&u(��wW�JX�dN�T-#�n��U��4\F�����#�n����l�r�8���iE,��wV�B�EP1�L�K��kx�W�[I�6�Q6K\�rUpl�E?���.R'.�u���ϱ�⽷z�RC��Y��Y���ybR��ܴ���D~/e�����-'M~��
����� ����W��!�3EՐ�@��/)�9�;�&f�:���JWr�˫�5�d���#L�����E��l�Zu�J����t���HC�Ά�����W'��,��7�\�������Z��H���*�	�A�_-�_�u���<6���)@����I�j����;;�1��?f�c��'�aʑR�
�	ܥx+����Hέ��Z�n7�[�/��zVfq�(���s�\��v��n�?��fN��D��c?c!�ݵ�g[d��N�s��\��S;ǆDzMYA3��Y�YQ@Ӵ�^����9�X�?!���Ss���:�*МE��= v���d�Q�=ኞ��F������:T�Vկ~%���#���s^��l�����jH�֝p�����ڵ̔�2dUΐ��RpmU���ȅ2	���v��:�>�K���#��Y���iV9=g���_��SY6���,������?Ҵ�W���̃ŤHjBރ��-q��p�)�@��+�$*����>τ(��մ��bD�8!�4QI��΀|�M��'��Sj�:��اe��@�.<+S|XC�Ԏ����<PK�5�m�vقHe|r`��[����Ǟԋ;��mc�+� �sn9�Á&�������2q噔\,�^�T����;3���;�
'�V�t���.x�{�>�U����Ȗ-+�tO��#`���`�X���"u�
~�MFGSv*3�V��RMbXf��:�Ʉ�]�~�F�Vz���$���Wu��Ϭ�o�C:����Fc.[��_��z�}x�9y��̽S#�NDn��z��:FN_/�e�5��G�h9�Vt�Ȏd�2��x�� ;V�-$�zw��z�����y6D�y�,c��v2_�?�0�v��J��1��Î<�dgt�ࡋ����DH��Ӌ�@�{)<k�J�ۧ�4�!r*�sg7��ԯQ��M\��T��v�O�l�$���q~������n�?�~Z�2��7㛆�5�B
�/����T��z�2|��#�"<����#�LoT¾�1��q1[�8@x��w�/���"�,��Q�1D�;���L1K�$��q�'�Uۡ�������81���`%g;��X�h�w�|SG�D�J.�i���!
�N���P��?*�N ��C��1�K�/��d/X��wF���~?��o/qxy�ܳ�S���	b��/ts������@��;��/)x��3�������a���q�ʹ9�N9�����'4MS���<A���6K�H���������r��tI$�[_ ��ET�����������D"q�d�+�+L�=�)�@���q�b�DrrZ��ޝ�	�|��'��u��j�Y���!��mbw�{�#�fi� |4�kM�Q��f0���G���4E9L)n	{�6Z&(��,���WT�6�r���1$YdQ���#�����L��]Q��<��C�� ��=M�h�q2u�{4F�N���`��:��f�T�
p��`���<�Qm���A�0jj5I� �I4*�U&e�˓4pl�W�c���1ʎr]^8_��.0�~���Չ������q'���ڇ܋2@M�=E�0+��`�Z��:(�5i�*�\���Dh�hN��ѕR��E�A������uӵ�Պ��,� �������A1Kr�}�#/��\��:T�G�gӲGLMLS��:ɻ�&���U��s�3ߞ��] *�w'gi&�Yӱ4�穛��~�A~������_�f!'���ux{f�
���p������MT�� C�ZnM��x�
��Ge+;��yU�����(�I��s;�^V~�NsP��j�BfgCwK�+U�s�x�-�����؛?͑ʐ�lYJR�u���7�t�T)�����@WK�H��Ї{�Z���HeX$h^��-�h���8䅌�?D��fkZ5�E�Q�,�q$�&���=@�aa���:��R��C��zU�����j�l���N�����d���:��zӹ��k�mM��X1��Lm�(�h�1ʩKBǛ���"�l}��J �}ٜ1���N��)6�9�#�� #ǃ��n�I74�<n�ġ�L�\��'6I�:>�t;�$�R_�ӿ�V��㦮����Ʀ��������g�B�I�R��Uᛤ$b�?��wþW�tnw ;\��/x�y \J�%�M:�Aj�^����8�������k,�I�Fv T�α��^g��sf�H���_,7*��DK�������ݚI�]�N�+���A�y��������j�#�V�h��������]���==kd�ַE��J��-l������K1�	� Ҧ��r���<���u�����03��p4��O޹��CyG��W�_C��\y�?�
 ��a�	�JҜ*�Y�Q�iuÚ���US끧�P$36�(����w[pA�[*CŔ�sth��B��nl�6a剶I)��}O)�J1�1�w���b6�(�GL���ȅ�o�v�9�`�;��#�P��g�H�9ٮ[����b׎7��+�GT���]de0�p�5�]��X�N^��� *��J8��k]�$D�)Y��!4��9]�NK�0k����4��O��'���q�-f�C�m�}�8��ns�w�yk�%}�ݯ�]�Zk�y��Q����Xk2.K�j���^��*�b�d �ޞi�y�?4Њ��4��LBR�(]�����K�0�����h��b��0Ȩ�k��K����%~+�GM�q����ɥ�,������q��'R�J�-�"|�����|�	!n��2�RZ{�@F�6l�r�{R�3��6s\���uCp���C�{_O��GlX�?���̍���? �>��)�*Xܱ�}�٪������b�r\Uo|ȟE,K*dg����6"~Z��?h+�EhwɽHt5׏����`R#X?k0,��|@e�Ǹ� �Fʺ:��>W*�𩌓^Kl]m�J��U4 j\�����em�M�	���Ӽ}}��T��f�E��&VAi�L�����ڹ�f��hz�+�&t�X�ӸS翃1�S��Y�� �~IB"�y���*��hD$�m�������#�?Uq�A�1U�&��1�����7��*^Q\�$�率&�	)e7�t�ؖF��s�v��2ۦ��=tt�'�+�:�F���b���DE�*K	�Z�Kuk:��J��6�����'Km�}xp��B�;ek6Q?�ND���ſ���'�%5XF�Y�Z�Y6����Q����v=,m�(������+��s�/ơc�"�e��3�����x�i�g�GP�I��3g�>��7~.���'U�f�
Ӕ��c��t�!+[�s���7ag��*CLg��̅y6��!\��\������Vq�Y������͂����a	x�赛D�|���O�qJoC@Q��Y��:��<'��hgך}���Q�#�ݜ�	��yo�M�L8:�c����	��7�g5�3�C�fOL���sc��<d%��0�z1��P�c?4�����/JJvS����M_���N0���T���7�^�&:Ev�"\1)���G ��,�����F�K��bi��3)�9�V�Rh�w��o=�r�e@xu27~�'��G/Ip���/�;�M$6Kw%�����I�O1�Xָ���0I(� ",\Dܭ"=԰�
"J��n��T�H�gtf��.7s�T��Yw|��f���=��f�=���1�7a�I�s�)�6��a3B,pNgk�n �{g#q��>$٘7�M�g^	�M`2��r�_�������XH!�+�̀�lj��b���$�iVC��\PΗ]��'�_C�~�UOJ�{_G8@)4��GC�S�Jq�(bf������İ
b\Q�*�y�x�l䅣	���jr����(fRp �	�N�]� ���H��;<^��?��'ϟt}���ǜ¬�>�R2�h2�Yַ�9����ç��a4��ɑѱ�Qׇmx�Ɵ*��c�(np;�,\���&R�v9`�ZY�2Ry��_i�'��䧲�`��n1��f"Ɋ�uI~�����s�=��?lX�@�t^�J���%#�O9k8�ǺLI�Q��v���͔���E��Q/&HQ�gӬ��/�DVS�Jo����eY:�!&f]	�V����BYn���zp��d�"��_8>���@QDf�,��Ί&��M.'w��En�O|��\�3ux�sZo}��$�+��E�(V��"�//W��޹/�}�Ì�
eN���Wә��l��`9���Y���I�Iz���{i&L�X�%"�b��7�m�f��Xv9���Y�6��V��W�][EF��;�P�i��lx�2/�i���S�؆������e�
.X?^x�I��rFuL"7t21�}�j_�jr���E8e ��T:���ߡ�8k ��u/Hp��5���м}�dH;X�������Ҟ��y�z��[	ؼ�:��&�>�} 鏎��u�Ek��M����rS��X��K��j-�qO�q��c�=̼o��Gआ�ׯ��e�i�_�lXF-8Ty�a=��W�[ �h��M�g>��U�����sjA��2L[�q�"�y7œXA��פ����uy�8�<=� 9��s)w�S�#��vLfgE9{K<P��$?i2P8�#s������J$v7L�	k<�n`t���������� Y��;`�f�n�TP8��t���1�૟�Ma���b��⵾BC���:=cHN�h�_D$6P�s�dP;�#/��4��%�CFh���*��?�%g@���K��4�.�d��pT	g�g��QŘ$�ڿ���@�;ka*���Mc����{:1����#A�K$p����!��wpI�I;"�_Tvqg�z��L9���+��%��[<�u�t���e7���rsCD�����%�� ��Z�	b��(�~�7B�F��Q�y���gv�ҷ_�����1��Z�ɂ�3R�|Pj��o|q�>�!�.T�+Ֆ z�?����KrF��td��p�>��w��q��k7pӦ_��8v�|���0=���OB��tL�^����\�N�ۨ�k������Pu�֋�ǎQJ���AQ_�.�B�F�PF�؋�+�Wg�֍ g���Q��S�냩�\�I,��VIk������Q� c�4`+X���m'\K�����ͬ�-5o��Sm��#d�yÊ{�Ǡo� "���{�����t����ш�ٹv���Jly���MR���-���
��ec������p%e� �j#�SX�~l,
ၢ��K��>�L���_������3�Q�#��1[��Q�*�e���h�C2���ڪ����ڜU���Zد�����_�ϓ	]s�_�i�E�Zeڡ_�q��'���V_]ÛlC�����`֦��5V�vP0�	��=���������=X3�����X�i:D��-�K���o��<.L���j����8�^��d������1��~{��*�.�2���^~[._&-��U�y	��fZ�ǽ�\��ѿ�m!�^�շ	���@X��-YB:f�'�`I����l�IQ�7T�9�۸��ȥJ�vh�nXW�z���lz_,a!DN��,�3FI���^��WNP��T��[�s�,�	��w�d`[hS�z���޿?�%ܲ�}.�a���z��o�T�l$T,�j:�^��A7�R��O�a�/��>���5R\[�$I��*�S��R¶�˙���;�~�1���&v�l*��A�q���5iE��(�g�����I��4���w2y0�3�	]t����ǳP8�� �osz�'z��fT��'F0m6iL��hۂr/�L ��d?&*̶sE�'#�yN�Q�M��R�I���H�H h�7[p{a~O� ��m�����<��IܟR�c3���1T�tm�e�x��[��U�7%���䯙�j�朙��cOzi�	��h-Sq���D,�5�wUb2iA���*��ci׍+CK�]>���#LjN�+#��������Z��#V�D�#%:��/� ��A�vxI��&R��l��`��֋TT��l鸅�`�0�L��)�fjE��g�=�*��w�Ƙ�a7F�O��m��^�㑺��e���\� ���	�zA��5���C�!M�h�})�װf8j��4+2�)��nk��������d�ц������jb��Amsu*r��c���H�$:��5��,�W|���m��@7)��=�'�Һg'�=�$\�i6.$sɽΖ�"�*�$8���SU�;�Dtל!Z���n����*�C��&�D����wR�����B��G�5�ђ��W��Ze� Q�9%���q���s�H�)��ˑ��q�!S��G%!T��8�JkǬ=�� ޠVUk���R��9��ClŞ�%��Q�f|�"c<���E�л�L�=5����m�/�?b�S�c�rj�ޒ@��%�Y�i��G����U��J�Qi��+�i�A�����5�V��e+Kr0բ0�P��ĺ.=����,��j��	h�?L���"I9L�C�z�|I|̈́,6�{�[�ц����τ�1�Y>��{Nz���O�3��iz)YP��o2��R�w
a����HDc|2����}7"�<x|�m�!�����Q3�5JtC��\K���?��]�hbVqL��ז��8#�Z��D]@	��B����<D���,[��}ȘX�?΋�Ȅ�?���,3�������9W��x\��q�bF���X����L���K��io��Ɓ��N���S�����/�z�0r��=��`��5��L��~��yFբ�Ulp�����\�WI�\�7�L��̈́�$�u�E��s�w���C�~���)xp!�B�R4���V���=�ё*w9$E~mz���!PO��ư�qɄL����̬��Q��"��;Lr�y:�����Q.�7��~𮯎ְ�!�.`F�� ��Q�U���j,�c�#�vj�򥵨 Y)���{���
���v+��J�ґX63�.u[8�@�vwKeJ��4_8(h���`a�ޮ�2ڿm��y�o2�S3���Wu��I]���x������*�.���y�}� с���n��-�8�#5w��=!V��R�v	�}�o��裎z0��Ħ�7Hޟz=����'��/�w�m��31�1_@�P�]��V7������	s�=+�8�i�v�C���C���>��<�������{x�r��	��A�Mz������}�%����G�F�8��f �o�#=D��S��X�pI#�rd6ɢ0��wO����K��\6��7P�7�"�"l��ӧ)��\��v�1?��Cp�IE��1�(Υ�5HM&�&�$ܼ�{���V�!Qa���c�S����
���Ï��x��W���AE*�+�e�5�2]
��X(�U�ᢲ(�b��u��x�8��g�B5�R���ħB��s������mt{k���jxc�Ib|���A%B��^��Kw#�b���	�P��"hͰ�[�5Y���U:)�G?�Im���7��f���_7��Jx����a�0�߷S�ԆO�E+� ���vLA�����ٰ�kO�V��Mo0��s�����N� �Z�4�t~8�k@����y6�������hT���5�LEo���Oސ=t[@G�8�t܅�u����i���>�#V��!�r�G �sS ��Z� S���}�t#о������b�8)׽s�����r3�0�xi�D-q��LՔ6ڿ�:��y>��t�3����A�W����e���d���NV�0�]�- -��t��%2�Mԍ��I�I��e����ns/g���2뷲��O��8��[+��ayw���Q��IKB~7
��8�h��M=E�/�m>�D�����w��8�.+�n〾�bX[�����%�a��*N�x ^�W�u}Q�l�Z����J-���tZ銢V�:O�5����P�	h&x��B�:�$��E9�0�^���2g��=�de��q�`�_���vf[op�,Z�%j5:�����7��_ǀi'[��hO��JY��o� ��it��q_H�.+o�Y�
�bŏ��0�ۺ��MY�giℊ���@A�w����L	���g@�*Љ�6�'����ة<�h�)K��z��g� ��/\���İ���'���`�/Ke�]�5.����ݴ:�W�9??��8�J:�Ͻt�}��F��׸��f_c�����/�֗�v�9i�����E>�ÜQv��8�1��^���d0C@w�S��2��l���ެ�������<���o�vU\7���Ik
w��hx���N|4�\^����ɚF��r�e"�4�R��;��F��R��#q��S������7���L2b�O�Ϊ1�޻�G�u�5�*#s������G(;1�y�A�"p�A�~^�=�O2�}}��84��#�47cV5�|��M[P�x��;z��	�a���	z�{h��d��	�*CJ�[��TU!Z��Ay��t��j]C�NDG,��4����$jBKR4;o�Ժ�`�KY��3���G�#��f���ݖ�7R3K�n��=�З0�e7�pY0�`�z�@%�$ h�=
 ��3��3h�^��
;I��Q��U��0�U�3vqDH�L^#���E7�@&�1����)�xtk�q=x�qAs%%`�
��¬y�m�}�il��&����\J�[d�|9ʉ��ʳ�y�y�8��ڌg̿8�^�[�<=T>$j��9�މ�"�Q� =�2w^#sI�5�&[q�CJ���:$�C� ����>:&�uz?>��cK5���Sy�]SI���F�"mY��"MvdDsMP�]������MD��I'WUvw>�#���F�F���t�q�Z�
Y��|j'_/S�+�����4k��SrN���Z��H?�=�/jw�oda�yIP��Jk�d��C�j��I@�����ш��7FE�'��5����x:1%sE� ��v�Z��7�n�K�僔f'�d�l���*Gw��^r�6f�0Wu��J S�ź@���^�bm�&� н�Z2H��rXʼ���#���J"C�`���.����J�3+�Z@���d���c6H,���̩��6�R��6h&~�fAo,G*�3��-�̴.,�x+\��wʾ^b�Ѵ��m"�K\ɝ�O��δkFe� ���ۀ�}|�;��g�����?2���qѭ.��6� �nʭi/?li�쓖ᓱx�ߒ�%�}�`�R����뎊���BQ�����DǶ��9������C3���&uN�;�ݸmb��w6��_��1>��m�M��萜��[@������Xp&c#��A
�J��{���s�A7U����e�I�-J`�f
���~]�_x�&����%�审����^�I���~u�Gןe�,k��c��L���Rс̂�E�܂���c��<�p���B�قӭ�Sh�f� �J�"w`_؀����3;꣹�SvWQޢ�\�4 T4Iydԟ��}��kP�\q��I�	��7�ˢp��T������R�SMJ��+�㞈d��ToQO����GXDZ������4�"ڃ�f�D�IS����.��]�#��qsœ��Nz��~�:�~z"tE�̥��奒����}�A^�\�+�a� O�[�G��0��^��a}4����ȧ(�GT���Η� ���V.Od�!E%3*M	{e�`z�Fp���>c�=�-�d-�_���/�x"�r��ZƦ}4�v��|�,�u�̜���4�&\��)L�J�~;GsޢsT�u"�N�c�Rn�S���h�U-��)�������I]_�������e�Y����G_m��h��Z�b>o�~�]�<��S���=�dv����"���q�_���!?��$�a�t��ĭt�zװ0��Ԃ� ��'hɲ��Ea(�V����2jӖϖ�Z�0QA��xX`�s��y-���͜����HC�#D6�^~����jU�='�b�y�vcR"^��/$��KR�{���x岑�Z��ǰU#��<�M��B3��y��Yl�n.#���U��B*��l�PO��J1�ڷ�c�ͦڳ���GU0����ۥ�a�[�2+�#½6]{�b�ߩ�� �*�Ǔtq���i��Nw�!m�E�M� yKEMG��l�/Lې-_n�'�Q�lMɫ\j)�Y�w�����5%����V�x!��#�&�|�ǐ��l����Q��x�m�ۇ�P}*ZWz�X��
R����gi��e193�xKL�����ٞ�u��Z���H]��fr���z/���ܘ�	xH}S0���ݔ>Z���X�u�{�ml�m���f@cM�9B�T��:A ��^1����!w�ȃ� Vš�����CN�m�?�e搾u�)h3Eܪݯ7)��g5w��s�;|���q���i�&�8�C}R�)�s�J�&U���U�$�W�"�B?.�զ$�ϟ�M��D)�͑���D� ֿb�>�mX��H��U�ŗ�ƹ���XR����3�oM@Z�K�����P����F!�o}fOw�L��4�J���.��1�h�}�g�� �C��7a�Ԇ�e�s�*�q��>8�V컉��S��n�8/�������w��3j�M�5�]��(u:H,�NE:�������\ƙ"�|�h��_Ҁ��^iT�B�'�wge��e �kTew�K�+�&�a�;���-?k�8�6���T�k[Z�ĥ���QM�6z��si��Бn��#~�kg����?d����4f�ak��>�Q�~�yp����{%]�2KlM���L��2��4��'�� W2ie�q�9oS\^���b�79h�٣D�)�x��7�kgÞ�}f�y�� F��!�"8�����JB����f�'�7��*%"�.�X������$�����@�3䉗��/2	d�Y�#�خ��M|sWf���.u�Z1V��,9,�Ggu~Y6H����~���&�L���
��!K��b�No�#d���Y�"u�5{,���K���(���P2;��� 6>�8E�����|�n�}#���.�0��P��k�����H�����G�� @D�����ÉG<p"	�Ƕ9Ԇ^%�0���R\���9�qT��d ����ǍI(�Bp��PE��4��vB$K֘*�F	��e���Y���=�6�����y��@U"%�|w�sV�#����|x9p��W&Yl�fCN�q�74��[x�ħw�_�%�ǰ��洆�Mhy��o�>@3L�ذ����#��p.U�7�M�X�J%
�1����i L]����͓e��<J�R���V
��9�C��zu��\�r :MV����ݎ�y��7!�ryo�>Ơ��-Dۛg�E�"{de�be.&	d��WG���&<K�r��B'NѣPz�2�6	�^�n��#ƉCY�*�&�ec�56��`Y��׌�Q�|��R�!���zS�[cx��7�5��n�5/`Lz���q�ͪvT�L��ͬ9�6��"���Er��{k����o��uu�\R>k���H�Ko �-���	��z����?-�X+� ��ilq2�)�1��YaJh�C3d�{��JnL�m�H�W$	]T��ա3WS|�F�#YfZza��`?�i����)S��$nz�)��ar�ib��.��0�5��J�_|�֒w;D�D>Y^�4�F�t����`L佺�B�w�G���.��!��n;pշ7�Y�W�"�����"\�攆�ÔyH�"o?�����W&L�^�R��(�k-A"2!�&w���_�.qRS�WF�U��FĘ_����M�9��lQt��1���F��Ƅ�<`����
gL� �*�@ukM\F	��(5պ�\�*�),hG͠{�ZTv�G�����J����mQ%*c�O`�RY�y��7���e.�:�B��܋C�}'	�8�F��8&��h�"�OL���A~�8ɣ�?��ޫ� �6���q?����e��F�����bR*��]GJ��.�!%7	]ʅa�,� 2���v�w�W��=d�y��Q���o�h���"y
�w�B�r%���T0�O:/}n��3h�4�)SR���Y���#��O;�
]�Ǹæ��'�=�0�Z��.x.�@���������:�B2����6a9����s$�!Ҧ�І]L����$#|*<�g���q�Nsۥ|ɶ���pQ�S7-�8Z�L��z�e�o���@�E�� �-��ښ"a>#Qe��'�m��4M:�4���� %K3|��|s65kh�	))������2/�� ��,3gƤ���άK�h��axkU��8����Y]~%��Oe� �����:���ҁ�^8�:�	�#���D_J������Xr�={���(��U�|8�F���:=����JƗp����p�cU�~�`�?6�z׫��z�,�/I<������J����z��0�ކ� �cӒ�7���$tU����i�({��{��d���̜*@h�J�����x�c2;����+N���L��a��dSҜ�������'3���U׉�:�$m��E�wBA&�9O�KUT��Z�.�0�F���L�"�5v⋟v�l��UtS��Խ�ܣ��J�o��3��{f:E�1����*Ȳ0�"s���f y.����9�A$d��y��}�u�Ƅ�^t���~S/Ap^F��<�R|����3�[O4	ι/b^��rƅ��N��:��F��"�{�7ӝ;R��ɛ�!nw�T���v`�YO�����
y5�i'��?�0��xpEU�R���Ie��X>y�i�ZgLK�:9�2ͮ�rp4�5���x�t�z!��#����Zg��Q�(Fx9=2��v�>�e��#�"��U�ĕ{H/��rw����>���EbŎ&u�z�s��m(�B��FO��¡�(�����ͱkmEoٱ�4&��߼�Nn.N@$�:W�>�D����V�A��~�!���=��)�`��LɲǮ2s�HaH尓y�MM����Y�W�����M���ϓG9V���,n
�NK���w��]k�|)�uR��}H{+_�vlj^�DN�≢c����^�:G�gk�~���ܳ��{1��X$l�����W3����?�C}��M�����Rʄ3t�G��7p7��g;��b�M�H�E���t�֘�b^(��K�L�	��7�9B��X�5}�|�_�Ce���&_?ͥ������'K;�^�-���G4"���[/��#�+�x�^�һ�8̭e���d�z-����,�+��@���Z�^�KU_�_��x�r:�Ⓦx��=_tJ���^֐U��3*K	�>$�8����KH��Z~Y2�r�<v��5�eN*&F�����9|�B���(<�7y��3��Y9��1��TD-;@���*��آһf�����зUx�����G�1a��ǧ Ĵ��5�`���AT��4��FFWt�]�9q�,-.�FG?ՑvBBk*�����p�40��)KK)��R�Eb�
&�Iޗy�UX���l��鯼ϡXG��o�۝0�o|ּ
WD��ue�6�vދ�2�5�͟��D.��=gy�%JR�׋��VL�e�p_�EғF�Dc���������g�\B��!e�����OP �=�?�1]1��,9s�q6.�|�@M~�6�,�D����q �^W��s���}�ktdZ�q��i�	Ǥo�@�D��*x��&|F��}�������ր���Ջ�	��HI!��Q��n���W_so�m��f��Q�C�2e;Q�׎��L�W�P�:�H��S8H5yE�)�:qs��1"����piv	�K�)��Ȣ�{��q*�C�Ȳ�e؈t��*�r$8eb�<@c(İFv��E=�x��9v���'�',f���v����A$sӉ�e
m���ۚ�)��g��0��S�@�c6���~$P7�dT�|Q

���X�Ln�P(�>$�p���$���>0N˒h��#
�*��Iu�`��a�(Z��lj��}N�@~8���pM�ۥ};��4;�\ɢ�%M�0o!?����@�TE��1���J���rȎ��.���wy��γ�X��Nj���S{�Y�L�E��b8�i�Gڂm�ڡ	.���k	�9~�i�g�G���*�����t�0,̡��]��(�7/Ƽ\���y$`ȝ�ט���C�#W|��׾5�DM�=i�@���%B*�8Cs���'-��Bmc�b�(]l�<����x�&|W�#����Y�HL9H8||��;0��������J�[�s;�宼�JI'�/R�x7B4֥�m�c��댆4�x�\�=���i "���m*Gk�c~�=�@��^��ɚ�aJ8D#����)�s�Z����z��#�S���Y��qP]Z4՝�$�:&���y����g�-�Q�����4y}g̹aj��	�Y�2yc��	U��z�X��c��dy0�߆�;$3+[v�L`���[��qD1���J�pB�O�w��6* RP�� �˥s͝�6��\�IF!�itw����,��U�:�L-V�� 	�~��N빺������ƛ��\����DPqJ� )p�tk�p�J_)J�8|G�ˮ���lX#c�P�Ӎ#�1my�SԈ��z	|,��t�']W���Q����3O��
��((�8]#[3���$�<�Fu�v���uY<���HA��6=,`��b@Îꊠ�C���j\�􋫲�=����Z��yE�gI�ђY>����[͎Y<A���e���)G�ej8��/�f�#���O��3�P��3k9��b��)ǣ对�P��E@��%��"�I���	��IY���T�#�[]p~R�~�	+J��MZ'5���p�yI�B��C0� ��YF*ǻ�R��bD\d:f+X��}��h` ��`���sݳ�������exC��F�ƭ��^5{�ꌪ`u8E�ܙ�O	�j�թ�8���ע��B>��r������կ���kȋ��"�vR7�Z*�aSc�<�7�6�n�1�f��'�&z�T:\���͆1r�w���=�V� ��H��b��E��"�Co�%עi�Y;��T-�l�����ܐ�vOX��	�y�Jg��2�_��{u����&��Z��\&�^�����z/�ߝm����v�Uޏ���?�b�I��X����"��m�����w�4���xқTeA@�L{���`G��g]����M�4c��t�sb�4f��>Q��#u����h���w|�(>�Z�k��k"8x�Bt� �Q-�y�)ػ��+ˀ��;X�o`��fn-���Oc�'s(^[��y��:�	��p�l�\��7v�n�"�U��e��7gƝ��;w��T����`mx���9��v�(���FN3���Xd���%HQ�������y��-EE���>�RYF�,k=�(ӛJ���j�Ov�yӽ1믭��ډ�k�C�r>k���k��J�n)���~���T��#%.�X�g�>+_-��� �����!�?����נ��S�]��I�u�ާ�G���~G}��S��	[���'h&g��`\ ,�'�TʪOq���T2���1��ȱ�>{�\�uEj9n�4��쉳�"��4�J�#�&צ��f~�U?E�z���n�z����g0�_{t��qϪ�"+�Z7�5 �?����5�Fr��U�|lbZD����mQT�;��%Ok�"���g�ށ/*�-]Z�\��8>��Hy��A�d��e�Zc]�>
č���|Ǐ=�����9���a�F�~��E��t�� ����/
� e��U�Sp�K42��U\�"$���44�p�#O�魈��C+/��N�V�4@�"��ϋ6��%qqp����9���=}zy�w� z��^�`�
۔|���6�1��!6�\
9�{��ܒ�`�L��Om�ɽ��l:����T�>w'�����#u]^S�Ϋkr�=���O�$Os��ؐ����H(�W�r���M�𥌈{���4N�Y�A�.����٬�4vs���$K��|Nx �u/����aI,S���I�o�V/�1E'q9a�K܎���u�%�U ��Tn��'3c�&���dS�YRPr����x���GU����4��8HI��ȴd��ݮ�P^���	:�2k]dB.�JGB�x��j��Cp�~����T��#FzF:��`s*܋����^� ����������T��E�k��u�>�Yߙ2�Z�����~��Q�5� ބ�&��۷��XQm�J�ƾ;�(͊���)hftx#�1���1f���;�6��H�y@�3i�9��)�.���Ģ:nҦ�f��1�+�@h��7�%fB'�X��NGɻc%9������miЀ`�ɤێ����B��&�#�g�MSW�s����@�v��,7O��/����)�h��mX�,�(�^����ja�;<�K�;֏'��DOnw��o��C5SG�f%jc��B����c�|^ptk�������5o�CG�V���Ҁi�rT!�Ȱ�=-���ﮑ���zj*Ɵ��1�-�YR�h>f�������4 v/*����6*�����-�6R�M
��#��uy�֭��$h$���Zo�y3�L}�׹UN�؀n��H2�ͷ9�~���7Bĺ����c6�}��V�Va�K����%޴Er ���㷆�7�M�ʻ�&e�az�����o�@��W赉��(d���&�ķ�!�d@�U��5|�e�)T3OeέV��2t�m�N�7�����LB"R|ğY�@��5��Mvcq�Cη?�+�<��반��6�碥���k��f�4�b�������ž1Y�_�Sa<��S��Ld��@EY�a���.�Coj���z�����̚��A2�# "��\�\-�)��&.d1o���f{�j����A�B�e��Rl�����f� ���ϋ\@�{N,c��1i�
��}V89��XO��~�I���x�Mמ�B��=����|thjF�5��$Oês�rf�	1z��a�i:u�a�EɈ�,�ם_���q��)l�b	V/	��(f�d�u�N�[O�#���6)s�3�JS�=����[� ���<�)�~`�EK�wG(�:��XϿ�6"(����7��r�ᚶ�c&�v~����!�U�>��/!��E�cr1~p���U�4	�#�S�㌱$[�]b���&��o'�Q�D�$_�7�8����͈k]w��a�}��I�����V�e`�!T\r��4|JJ;YmP�>�?���,�SB��*}�j� ��_9�ؑ\�طl+���H/�:,d�7�w����@G
��âx������KS�<��͜��{æ\2/D�,�s ��;2oQݣP�ǯj_��X��r�ڬA�M��s���}�`�xB���+�:���&V����2���0ld\ͬ�JZ��s�8��*��S1�X���	�� W�NX��V:����`�1��TAt���{��U8�����a�$�R��%]�����3:��ޣ�������i�0tC�љkԭf�89	��KxU��+�w�Y��`�������K"
�7�~���k䧃<ñh�����"k_+\g��<�oCG�0�_�x�W�H��2��c�t��G�O���g��wSe��iLZr�wZ�r��2��݀q�1��+6��̚@~;�������O�qyx|,�&�x���5Ò���Rno�6(_}�S��N_�Ҷ�Ș��Im���;�~"Ν���t5L|�VBT��s]��́�_�����׽�E(�H,��&&҂Q+'N	��B��z���iw~��NϠ=�z��Q�p+]�m��k8Q�&�b_�L}���WG��IH�������yF����Sa��B��1�O\ɜ��8?��S�Nf��zea�N���#v��UFۢ���tX��mwY�]j	bm��T}p'X��́5k(�UBl�9�!�T�W��mb60Pq�ѿ�F����y����O)��g���wڳ���J��'�%����#��M����7PB�O�Լg���r�v�_Ji��>uO?���.���rh�o���nv���+О^�la��t ����qB�>��h�h��z\N(����
�WWG�k{Ħ�&)8TC�l�v�i��}m	x-���0J��q�֯zr)(�e���2��0�M���6�ú�m-XwH�x&����t>��-e;���� Y~e߉��L�K�y�He��J��ñ��&�B���H�z5zOU���uk5|�j��>{#z�|��\TL�!L�!^[�-�E��Եl��?J��I���8�}g�G�yT&�w�&��5iu �	lyY6������*�j4rG6&�_�6Ef��e�x���a����2�U+C�����K(���p�����⫃2�PK��ɼ�U�hgU�Hi\���&�2�RK\�{7�.Q��{��%�
��ו�rRjн���䚲x(��Daz]5�*�u�),�2,9�0����b�B��XNx���`�!�V��� �m��/�mU�Ӳ��x��<l�v!��2�*��j$̦5e~�9�}w�er�n��\���@����$5M�M�u(��:�[���x'Gޏ�Sb��2�/t�v�P��I�'A��sd�hdr�y�.Y%��xBN3s������׋��IП�(���_R',C��B\�6A�ZMQ�n���ı,�u=�f�,��r�����$�qY럏�1�>�Xb]�+��A��@��,!�s� ��F)빠U�|וg*,��ĩY��p3�e�腀�K7&���w:�|:C��x
[MC�
�zwT���������tl/vz�����-�3-I�Bm�t��s��g?���ey�u|B)��4q�3Ypw=0b���K�p՛C!�)��Ӗ�4� �I�?5^z�Hn�l�oZzc��zHmJ�oc#�������M-�}��uU��)ub�N+5%��][�h�Zؓ�-�Dv�P:��O��%��R}�J|x�->-`t,����!�LU.\�H��m��;H��X�.���7Zm��� �)y $�E�R�\�=��5 A�cQ{��c�����ZX�bv͚9:E�.;e� s��p�2�c��_��B,u�bu���$�cl���TW�ll�C ���-�޽Ms�Y�E��g��&�bv7ܡd$���e�	�;��{���hY�1o���q?s.j"b�Q��\v>HJ��Ԧ�~�$���lK&�EߓP�7���
�dmʫ����Z���*θ#����x�2��w@�� �
M��lܣ��}]���|�>��'�=K�m#���EG��n�W�d�{������=��S���X��c��������i��f����n�g���1j"q�)9���;:�}����y�c���a@^�*x������u�����	�\�%3��՛n���(1�lo]�c����:;�GclLxb8�����v��b��"ɹ��=z��Y*�!�-B}+�Q֬h+0e65e���� ���}�O��tmh!�{�aN�%B^O�i��]km���᥃/�nݵm���X05�ϝ����n������C*Q&R�Y�aڰ�&��\��
gG�����%NsPn'�=J�V��'�t豠[�Z�����a�1z칻��j��X���bWO%�R@x51��'Ԋš�9Q�ʻ�� R�笨�#K�'a&�dʀ�2�%�N���ɶ�)��,���rV,^z�|4�oq�=T������o�B~eX��"�N<�Z�i�l�Q��]N������A8/�g�,�,0�1�� ��03�v�&�r��1�e���%�l~���ϻtg%w�X5���#j�Ⱥ`=JQzg|$��գ���G\�����x���%���)Dm��������L9#M����WI|>r��2�̻���f�;��g>��b�6E�pԎnַ��W����γ0��(��$�Q��T���P���1vI#J��@h�N�7:��p�����I��&s}2xY:%�ǀt�^m<��ܲ����_���.�xrT�B�4�������s#���y��y�<]SD$���k"��.�m
�� �))v�DvqN_���s�w(�/_*|i7�pR �Ցi��|�/��8U�9r�U_���{�lB��nړ��6#��H9�蔍U��Y��k�=��%�$�	�u\��:�\9%q\��$� �Tp�ޝ��e�f��W�c��	#l���m�a�����N��G����i3Sl���z�g(J]��S���ѭ����fC1m��oY��_#�"���������_�ho��{E��T�#&d\��[FYշ�׽4l,�j�D���Lȉ݀��z����AI�F%����J��C��Ntv���$O�s��}�0���H�rn?�fִ��f8����?�q�]�^�F}��#2��p�	�����x�W	�_m�ܚ�u��/����5-�ݲ;)�*b}��Gn�u	���[?�.�{^٬-h�2,�u�e��]Kp.~	�͂u�����F{Si8��y��˨--ڼ`���"3���(�C�9�l�u�%���Q�~,
MaK��YC#���c��=��y��^ �V�S�c���ڣx�p�T����1�\n;Y���c�Cj����_���ῢJ�5���zK�]
R�3~,�ʿ~U���]-ç���hV�B����F?�N���`�ɺG6Z�l��v�"�D��?Ц|��1��Vq�&SZ��_gP�����.�c��F�[DD�3�^�Y'�C*ρ_2% =n��0c�Ϫ��leotzvr���j[�%,|B�M(��b��1T�ۛz�2e��噜A4��˙��(�R��k@ >���ڣ�_����i���؀�k���Y�����"c4P'�R�!}G������%�Þ��\�&j���b�����t��!Z��"�g�0�G1� �%l/�}�f��?%8H| (��Qt���j���%O�P�a��,^�cM�$��5�L��eC	��K�%Ǡ�WRk3�U��7g>�EO�U}ɒ�_C�ω&�H��|���י����*�m1h��\�����B:٩�~,�#�W��+xĞ ��+�ĻF>𤋮��	�M<�%_;������":��G��u��'�kb�z&�M�9�A��I�O����5��G�*l���6��-j��y���4����|��sߨ�o^����Kb����q�K�!��??m�z ������WdS�w8s����L#'Yc譾Y� zR�ПV�4O�����^'��	�b�h�������3���D�W[���F
�W�v�䚴��Ӌkb�uچaq��ɉ��Z��H�U[�Ur�gY��j��BI�ˠ��杪?��7:{�)�X��ʙRK��eܓm����Y���{�6��c��5��^�C�*����h�ɍ�N�b���s�FA���$��x�]�rUT�.�����2�����@6�O�c5o�Sm%	}�j�aR�c�݂��:��dE�>v#!D#Q��[Nb)�;����y�R�<��Ҕ��"�L�a���� �P0Q���]���^�ҿ��"� _ӨN��nK5������R2 
k�Яo���np��� 4�S�h�͖�ᾘ>eõL*��w�%�Ykl����:� ��׭!��A:���䱒�,LW�HN]�1��Ď�������z!�Q��5��os��-���PR*�NZ���:ǀ���?~S`u�2;ǪvpًR��QEȊ��¸�Y�2诂�i{�C�17�e��+8��0��q�e}��&Tr���CN꣸9��'i�h"�B9�#w��������^)O�XF�Y�W�u������̫�nѣ��YJ�׺GY�,t~rѲ�������r�x�@��C���	��D����>pPC %`|�����cm��җR���l�<�'�5e�j�v��ZX�����9��vRWx\|�k�C����@��j"�����o)�a��/"�T�@���5�S��7�Y��`�r
; B<F+{;&���7�QɼM���q�~�J'b��;��)��2b��"��(�aMB��7SJ��9�nv��J�e]�1��x|��W&�>�њA�_�0�m��4�d��bL��(hk�o���>��`���x��\+"�V��>6�Z�}`5�+�wR��]FP2vzْ�]ާ�4t.z���� �V�ˋ���b�DU��I��<����R��.�d}nKLh���.�������:ƵY��d�ނmx�ph`��q�N�x�������n���]/.��2YQ�&�؆%���M��%~�y}#���Ϧ	��5K)��+�nS"���Iy]��$��X{z���2�zxULD�J���6�Ӡ�x���e���S�7�w���4qt+*XL~�PK$�@�r	��\u���g$������a���m�A�ä�h�h�ܷ'��W�&x+nU�	���ċcd��Y�A6��T��T^��׾���!�@k�
��DqDM ���5G���KI+��ёe�|dZP���쥰#ͥwCW}.-`4��&�)�@�B09U�\� l�!(�%�"���u�8VA��",���5������醂���a��������&�;Or¦w]�k!t.�NR�U�_G��f��Ce���XJ��ow_��S�T�!yEJLk}+�i�-$>�W[	��F:.�Z�Dw���zpR�.�Ŷ�L�p��l�{HM�ݮ(ڕu�.I��:uO�5?u��-�f��=�C�MG�-
�)��4���^�;er6�8���b��(�S��
��e�t�z�I������G�7WN�ǎs�'�z���)�"�>@Uk<ЙF{^x}&k(��'_%�%�+���t-Dj'3.�)�dB�e�����s|ت����`���i��9TD��dF���V^��p��/�hǗђ6���:��8� '��/q��O�	�6�Ά���ik�3�=����W�����|���8	;���a�����}�
br���x�P�v�q$p��̊
4�|�Bf�+ �п��}��(�H<Lu�6��h��_Unf��7��(/HG���Ϗ;5C���P�u��9�D��C?���#�#_�r�a�YT�f�ًF���8�Ht}���\� [Z�^�Zn��$z���r��uCH_�k,�Z��,�7���`��p�K�f�'��2���{x�o�x�bo�b�@��+~��m�j'�E,mg<t�p�W5�}��������1o}��1�FT�n�:K��DM
�}�������-k�~d�>پ�?\O�Lz)�'{�V~�w��H0�DH��+�X-P,M��m�ZԜׄ]�z����VW
X�Gxv0��ڕ��Nx/W(�f�E�b;>v�*г��� �#f�<h�9�y�-�	��~&P�Ǉڀ�~xa���Y��V4j{G�����-����q���j�Ĉ�	�xrN�"�m �5��9�<��Hqz���by����2�T���^�ӱV$��h��e�g���sCΘ<���@J��G��_?��K�^>{V���X��Еn@Ќ���En��؜�o��9��y)�r]�J�/�3��h>�����@u�ՌwY1E�x����*�͂ȏ��Ȩ�:��)�S�8�)�Z��@\08͇�C��W����*��]�V���}|�cT�a�rK5��8Ғ#0�!,�#�����ƈ�̱�!��\<�2S ���_��K�Fn_�U��3~_����q�W%J�3��9�(�w��L��w�,�IoA�C�����f�V�.n���7���	��w�o�g#9�)� -�������M��X��"T�yLlw�7n~�{?_�s�Cz6c�;�<B�9�n�m����*��r��⺘�� ���&��k����G�P����˟�(�!�7EQ���7*�W$S�ekC���D�~o.ik#f�ݹ
��1��/MF���۩�M�T�0��QlO�H�*��}��R)���O<�Pi�0��w�:��u�9߫xB���C�����2�]:�����1����l<�߀�2鹑0-� �c���\�ղ�n�QMc��lϼ��PG��I��J[\~��,�j�ACn�q��bd�u��X���ډ`Ié�C�K��ɓuWH����+4�RX��{��P-��}��$�y�|�C��v�f0�NG_���~�ɂ��R���Yh�n\�	��*�����#����fb�����E R1����6��
�K�V�0�[j�iJZ8���f�+��ZH�zl.n�E���NG��
�i<r��k�_߫�8�[���nX�W��(k��燢�P��*,9��)E�\����=�g�J���BQϦ&����j�	e\������ڂ��?¥�m|����3?Wċܴ��xqL�,���9�"+Nõz�s����s���UP|��$��~R�&�;�\6� ��$UR�t ����)�N
4���NFz�Z؋9�Fl�-"G�~C�������#7:��R��+fX�ȇ� ��-������ަ�fqx�R0%�.�"Ƙ��h{#�^З5��!pC��&��ӏ>�KED8iv��v�'�����[�4�h �r��=���^�u�����[nj�
e��=��RyN̒P���M�L��'mMp?������18�/$��A�x�X�TY�W��;���	|�����u��Ṵ���aJX@
��Lk�w�Y{��A �M��W���tb+;�t��Z�,����?�d�+d����j�D1�;rR�+�p]��hL193���7�GD}ҩ���J�=2�E3��b���ҏ�3�L#f�PCZ���Μ"I������{��|���C*Q.X�rv��Q�Ԝ7[ʕ<��҅ xi��h��������7#��3�
R���P���f�nt���n�x���9,�v��6�E�ݱ�?^�e�]��$s��"��c(� @�;n&zN���/f���Y ��"�����3�%����QР�l��B*�w;%� ^������K8T���c��;�� �c�)s�����ŀ�L�#�L��fJn.�]�-ؔ�Z��/�_�Y$��%���������B�U��%��ע C[�+����o;��R{�A���R1�T%���t'h�tӏ��gx����2��xq$�a��&�
.�:�z�;�',�"�Z/	��n����˟�ZW��"F� �$��	6�׼Q~I�S6D�D;�5M��vk��.J�`�P���$��Z�U�t�y�V�1?9��uñ�u'�K���S]<eS���mvMA��m�Z��ƫ�[��e:�׶��|�4�~��9�T�{c1���Ac��h�摢�'+;�N����3��~�ϺI���C��:HO��XALa�6�]]�l\�X}��V�,�:q6\�3TEr��:&+4�,�oU[��,�Ei�8I3�^Ps��	+��9أI$n�����>�E�UX�o�Y��&�\�w�3��Ѧ�&h��}^D˓����$pK���%Iǚi�d��2 r	�Jx?t4�drT�#�0��������CT�%����J��d��c�.��i�^��"��ܞ�cδ�?�p�LH\�z�/-c3+R���s!y��p�~�?O�&�־"^djz��Di8���U����,����O�!�DO�<����5yjj��'�fp���O�F���#�R�:�1y��պ[�Y,�j�D1��qb��[P�Anq��* ������<A��0#��@����� W���Y�h%4�ۭ6�펲��@�F:���8�	���D�35�8^Ԏ�; �(���@�/��8 0�}� }�Z����������'ɹ�I�����hC(�E\|pu�,%f�j�	�{�6���J���8$?J����h���m5���Ex���v�����o��4�$unPmL����hG�����N�;6/@W�7��h�G�`�_��*�����p��e܌'�Z�]K�e�?/1ˑX�R���0�[0F\O<=�Y?�����0��.I��
ey�ⰴ�b9����C�t�Gi�#|K����LV^ߢ)�ã�G��D-�0�5<�ژ.��N�i��Ѯ�<��B�w��Y���Ks|(um�i�p|R� ����n���Q�9N��_��;�6^�6��L|��B��<h���`ڕ��h���6�A��� ᆮ0�e̼���xK�a���B�-�h)Ƨy��Ӹ���b��*2Ĝd����3��oDC$�Ĩ4O���3�S�IW�E�]�����-Q�a�8i<n���{2����˄�|��au?펁6d����s��B��`�x�Ӑ�q�uA�3��/�C�A��l<�Da/X��K<?�D�fPW�T� ���8�l�Wժ�w�)s4�KQ���K��>W��WD���~b)c�a�r��[�!��Q���-&�īNf�IC�'� X����^8Z	꣺ }����|���j��J�rhY@$T�D��A>T��R0.�5W�ڌƝ�����J��A��I�~��37�R�;�������C;y̭ ���)��i_�� WtPJ-�Jj�fH���k�eӮ[G���S�:B��=����)S�ɩ�b��JQrqJE]V�"���W4 ����\wR���s
񦮒"���J�&M"��MðHD~@���-�r�g$��F����\��nC�ܽ�-R���L��yGޟdW�,�$������6��u��������`�-/N�-�=~�dƶ��g�5*ty�����Y����xy�=��R�W05�����+����Q׊wRB[��%��&x�V[�s��T�z?d�E&�e���X##�,��;Q�=8�J"u��δ�Q��g�?��k5��#��/0:H$����<�<|��I�݋=t��u�צа}��.����Ne@wE"��ν�ɾ�\�?)Lސ�[����Dz���S=�'�+ɵ���Y�8��^�5�ZO����q�[�n܌)�����H���i`U�%�w�d	�-h;�X�/������q|�,|A�>ޖ�S��[�Cc�A�g|����_'h�\�>�����Os�XߨVe@J�;�_�=_)���_�}�L�4+��ҭ�|��mI6`�X���H{�w�%�c:LL׫aDR?i�>T���)��i��]g�s��Q�$Y5��A�۔���������܍M�΂��W�О�Q��R��|khij`�k�@��:`b�q��7�g�e����Ag8���s�1�Cwk"j�
4&��#OY����#���ˋ��'<6�h�>�K�����7��V�#�n~���%Ҩ�K���m�,s)�&ǯyj.p����o��dM��ɲ��*�]ͼxU�o�� t�z��qH�W-B|
�I�����ϱ¸�R}1=ƥ�1�{|��z���%�-X�7�	GP=%2o��ł|�{��5�<��Ȕ�o,��bW����VNb����l������9UO�H�"I������wW����������QG�+G��>��gN���}�����$�~�`L���z��o��O!%W!�ń�6<��	���`7ڿ%
�`���@�ZQ�$�_$e���WK�g0C�/&���d��G/����=��طQ������7jİ�,z-EI�h����L#@*��U����*+�&����hB�E+���Ye<�ѡi�A����HIJ��y��Rܗ��^����+��H0{�e *���
J�"Jh洣�uV��o� ���ߝ�b�T��$��=����!���������ޔ�>�W_~]��p�)��q6�M���-�<�TFȄۇ�!���蜗Fɫ�$��et�k���GP���e��d�&��yr��v�m[C��Y�خv.�]mzt����p�w�_��s͛*D������\�Lt$o���߽��!����i*�Sݴ�Š��ѩ��!���yRT8��x����;6w��\^��ZGN��q�G�� ���U�k�~0����4��V�4o��B��C��ѥ܁��c�x�OL���}��K����{��tV����7�ȭW�*j�?o�*�6h�X%�,N��%du%F!&�161T7"c�b��O�Uڳo��`�-�F��̣����0Y��R�V�DW���N޳���.m���\tN�ͬ尷�aqo~�v��qv���)6����1�a$f��6��Xe��1�^Q��FF����
E1d�:N�)�ooP_"4Ǚں4By�� ���"�����h��'����LiS~��d,V7Q=b���{�o��w�Wo�J�{ɕ���A�e	�o�k}�	_���-Y�O�^xz���������=)�_�mء�����[/��툍�Fe�!U?��==h��� ��s����"���p�_�B;u���w!�)֜R�
���4���V
Pu*-R?+�9�Q_�ae��|89X�+��������g�6cK�M�b��Vo?����{n�u8�ejD�=N�mS�KE�H�ss� ����UA;\� �2�N���+t�ƨ;����W����E�'�-�`�䞲�8l܍ߪ5����s1#�mo���RJ��{�%(ͱ':�lK�E��Oc��n�)�%�����7+��9�/̵��[�ݤ��E�0�4�T/�e��S)"��0��eV�o�J2�z��N��ԕ�-~�����'vI2o:/�A-�K�Y� �o������Ti,�]�]���*�5r���Æ�<�Ҽ��G�-�����r�
/Q��[%-K�-�4�2��*.Qp�������]�1� Q:�Ap�^s�et\��l��+ރM"�b��T�$����]O&��735�=7�+q��;K U�@3w�?�d�x�k���|�5��W��E����\��̼G1�2&����V3U���Z7�%&�C�ϵm�Q�R��>ה)<��|�մ����~��V�}� [a�P��!LB����s���:�a�2�����y:�V&�˽P������ �i��?+�T!C��	��G}
vˁVB8*I~M������p=]XQ�X,���参���0V���ɟ^�7%ACJ��*�(^Z�Gz�?�s����3d�X�~)�x?^�r�R�q{��i�H��0x�@V�L�	jA۞/��>g��,:��s^\��L6i�/L&����>g �A��?�Q�̆���2��-��f�.@Y �� ��5�i�8�z����ɑ �/���6k!��5�7:R�H,��@R��HN���O"��NdB9["F�51���"(�t��!�$�=x_6<�ȺR�~��/�u�:!UqQ�)6��I�d@���)�8�!���[�9ǨB�E����N8�;bP�hC�誋ϗb9,"L�+�о���ݒ�eΞe�\|f�S�_�@��r6-�>�S��U��nrz�P$���O���u�
�-�d۳po��I��q��ۮ�@�֐b3ћ:vz��4���%����«�XzI �n��GL@~��x�s"�yd��{�0��F���5��$�:��a���w���	���
�_�����ް 3SqG�{"?���]0[��ȝ�l��tR�	L��>w�F���E�\�+�z�8y����&���ܤ�dV�R�nͱф�Q��"8�����{x�º4�����7Ϫ
~�V�N��Dy���/�6��1�v�?W��z%���1�As��bYQ=��̯�T#�6�k�}�[�&�k��p�K���o��Gk
`ߘ�X�lW�R���/�s���;ޝ�T�)6̪�4�`�yłL=�{883���څ����S�-CG�������ǹ:McsP-��?�^�n�oRu�z�;��K1H&s�2(D��r�C�e�~?�������VdI���vm� ����*�)�pP��q�~{��>�<���F/io�M���\P�I��d?he���u�W/+Gי8}�>��������6m� �ga+��(����V�6�΃����OG�+��sV�qL�Fҫ/���!�Y����}S?��ܠ	��#�vDK1�: �R`��*v�hr=yXk�̓q��%a6��L?z4-�;�����ju���U~����x����Mb��dٵ�C朣kWH�C ��dz*�|�n	���
 {����k�ȳ��T�푳�{Ņ�fپN��ђ���Y"��,�E��b?GLj~�4'ܠŶ����?����F�U�|V`����lL�Xﷂ�/=�c �~'�\A��E�Ђ������~3j���\���YӼ��J�������e�H>�1ҝ��Y�BA Qҫg/{���R�y���.O�G\zz����M�}�V�WT�^hA%�!�G��&�D���|�P��SA��Kґ��M3��JB�#nG�n�W&�O��5aO�+������FB8��$u
MJ���.#&��gdc` c HU����5d~�97��'>%���#a���&����j�2�6�����+��+������T0���̖��ٗ^�â�h+ D��[��2j�u�}39�1�}������J��.:KYNo�d5d���<k�|V�z���خ�=)J�2���y�޺�t@��#�NqF�i׸�䧖x��c�����k�5ثhv�ŴV��Z=0獟Hc�sBw{�1L�ǡK+rs"sL#8b�É���/?�&=f�ϘW\p�bX��l�UPEtYBnV"*�\j6�����$ �ɳG�� ����|�e=�<gn���uQ�0by6�F�[?�¤zΨ������x�cno���Q�Z�p�����s��v�ے���͎N���� ���t4I3��C+�$l���K�I�\�
fn�#���O��H����_��N��ZTY�]R�y�EC����Ն#$�I}-��6~|q̓�J8J��k��
N�^�ǉ&\�>*Y^w��^��_R�c��z2��kdb���Xno=L ԰.�L�)>ϟ+�a�@;���u"U��'U%C`q���{foCW�?m����2iZభ����9��g¸����}9�4(<i���i���e�;ؕ���712T�NF �,&�J�0��]��k��X/Ʋ2ǿ�i!����;���+���e��gԄ����?Nm3�� П���F�~$����<g`Ⱥ���/j�^Ӂ#\ʎ�a����n#��\��!M蝏8���B�5�"
�4�e�s3˔�Z�NP���z2r�-��-Z�盛{0�&�f0 �|晟�m��,&�m>نe`�z�{e����I���*粀 ��K�~��T�}-�F�Ua���#p�RU���*&i��ל|�MPbv���g�ֽ>�]�
�JL�B���<�ơP�J��j�>A�e�Z�m�w�sg��)Z'm@WcO�;�k�C��	��5��׻�p,b�BĞ�A�嘆Lq?���~�lj�g���d���\Y�r)`��DK��#^@⪾��b���/3n��.�������[�̄N��w���,�5�M#lAq��p�Hp�����G��X�c��!����tiO�g��6�^�����'���LMN��4��<���V��l�O}1�S���+*̂�Ge_��C
�t�g^ � �ڲ�J�c=W��)��//�{�1���&t/~d�@�˟P������7Ã�:����z�\���#��6N1���ɤ������8��)�R%�g�0��G�؋����1���)��� @�7����M�s�zJ�|A�&ͳ-�l�Z*kѮ�U��t;}7�̀�Y���DT�5�	}�4��;���J�XRsja� Gb�[$�==C���b�}l��S����4�i���>|HU�Q�n�Ӟ���9��X�Z\�r������^��xa�m�9�t-��"uMP�y
�8�#=�C/��[�l�<��ѷYU��b*�Sj��ې�n-'��`�ްg3B~�
�uu�:R���̝P'�Pq}s�+o�f��p=)��	�ݏ� ���s[|3�}�6i���i�?yݍ�5�9rޛ�4a��vd+��^>�3r?\%qj��<� �kW����od�{#^�� �*a�s'*m\=�F�?;t���f7����c��a"8y�Ǒ�]_�'W)�x�Uw�|5�����;�f^0�f@	��CG^����8����G�L���?A�/�b��R���^�K��q��y-���rۋ=�69�P��Y��9rW�Qˮ�lS�G�-�W+���W�W�ǮU���m*#
���}�*��=�K��h�d�vb�Ț�hR�ȸ=�n�	�|�ωb�|N?]�j�} \
E#��.� TJ�"or�M��L:{N�޲	���BBN"Q���t�{]z�vˀ^&:����v'\� �:�2�j[�9��t��������F^�	��R���v�UZ(�5�k�y���3K]w4��p>����l��Y9����L�ݚ���%�m��=C���`B	��йFE4`�R������Q*`);,|�֮�<�"�5�Yt^������	�V����7���q���b��ڻ��@��=	D2�<_�.���oԟc�+�I�m����Ǐ2���eG^�/���s�ycw�==�b�JDٽ7�=? %��2�Q�q�E�l�Qۏ��+=���=)L�a�~8M�#������c�g��7�5�D`ܲ~�~*{g�h~8\@��s�Y�Ks:�r�t�mT1�4i��@C xj�Ο!�U���1I6�5�p?����N�ˤWa�t���U~��q����}�KO|��7�="Gd�-<x�������X�nR͎"��Z>�㊡M����FX.���A*&��>��a�t�<�M -tynB�}��)�u>O�f����V"k3M��m�}��`���0^j���YS���k=f��w�3Hu���5?G��O�XU�s�b�����1,�P0;�B�SL�χ�"�ݑ��}V!����r����ͰjVBH\�B��\6P%Le!q&a2�D���a�BK�#�\�\�3�8Z��A���.'��m9}�M��/x�y-P�_�����_%(��2,�""?Mƒ��{1��m5�D�h�Q+�Cnt#rݙC{><�G�ȎЖxՏ0��A�*UW�n7��o�Jp����!h�ߘw���E���[ٿA��#��T�L �y&�]���ZK����n��������]�cI�Æ��j��_���x?�u����x���쳼�x�:P偑�^�{�n�4�3R���j��"���#�J�Z���KwnC�-p�c�m�ˮ��2�MJ�Ls$�eLEՠ.m�I-6s�xc���w���y����us�Y�8��	���/s=U�|�/��C������XV+s7���N/;�k���\@��A#]��ZkZT�FR�4��k��c	N\�QąՌLuf�J����}B!���E�:��w�^�k}������[��\,��)���>9R�5�
���"�u\VE"l=���*,��=/��M=t�D�A�>�}�H��S~i�+�)3��೔���߸}M�*5}���ۭjs����
��i��&�r U�D
M�ݏ��\ɜ�]Y�+���I�׉XZ�:ɩ� Z�)!��4�4C����o��As�_�j(�b�J�e�`=?�i�ciR[pOE��P|޶�>����j�J�IdD�.b@�D^{�˼xI�(��|��Z =���%`���S�;�x�$ș}:~�B48U7]���s���&հ�r%�P0��C�s%]3\9Cnl��X6�?á��L4����� Η�"/����w-,����YP���ܸ����g}�l�oq��bt׉6����: q�Cg������G�L�7Q��c��(b�`SN�b1�|c�:��\/?<&��9Sh��gY�ޑ!�{�/�4��e�O+�P�@���T���E톛N�KE�/5�?a��
�@��[2xS�=�q�k!YLT}'�˴�4kW��;�6MY�W �̳A�sB��e�ç��K���@J��.�#�m�%;���y��B����^�	#6�0@Џ��p���?̜��ʎ<�S���@��u�O���ϔM��oZ��)�Jr�c�����' ��>N�f����uH}�ALI�9"\{�k=}4z4ugn���D۠��e
{�Z�T�]jq=��R��{�}>j���E@�n�{�VO㛯�&vH���o��O_T��[�J\��$cxLÚ��M��6dM�e�ψQ��f��]�=d\�>Cj31��Ǖ��j��~.��=�m�w�n���~j2RƐ3Eh��zo��NG��v40r���a�$7Dܞ�����2��7��d5�^!��/k ��c�2�y�Oܜa�µK^d�,(�>�Q:�)���:����j��[iU�ŃfF�Y��4��\���?���� ���I7�ǚ+N鋧5m�+&4{�Q}�d�DI��d�F���̫���W�o�6EmM�ŷү�5'����tڨ.R��� !R�2�Yw}�Fu/��-^��r�*�;��Y��V��'���f�J%FS��B!T�q��:���?c���+"E�IET�7tk<�cc� 5�f��D�a�
���v�WSb��:i�RGM�=4� �,+ːC������A�)?>C�T��!�էp�B�mX�֥�~��0y(}�U4	��]B�IU�3TD<I�i�͒�+~�DMwJߖ����G��W��V����xg�K���y#K*1���di�U_��}��S5�X再�8O�aW$hR��
i�r�9l�W%#����q��+���d �#����Z���d������?x��<X�/"�j���YeG�IÀ�yV�TC�⑆��/`��g8�D����>Np�q+3�6��h�sg@�>3��9�kڀ*� ���\R\LG�֩?a��=2����m�����炱]Ԝ��ʋ��.K$ǿ�zsN�g6M%Y���R�c�7Ji� �~�
x��㤑�մZ�o �òw�x7 �V�� (a%��/0�*�I^QfOt)� ��ͰV��:�w�Âʹ3Y����7��{����������nw�b�D@\w��(����ҿ���%?dA�"୩>��
C\�Iɨ�i�A�ꅟ�w�'2�ڄ�U[t��U�A'���n꺍�e �GJJ��5�&�O�F?	.y�"�lY���Ar/aj��4^m��gmx5`/�W�n�g2I�2�꟔�K#��@ag�*�h1����(�.�� ,�E@�&�$����z�_䚇�-��P-���x4��p�e��gow���g��9�}�ۨDx�:J�\�Y��5͋�}Ф-�k�۰��[E?����;�QQ<�
�V��T0R��A��\"��vV����r2���^��ߣJ�݀�N���)�|�k}���/h�.�s��z��6�+�yA����<���O���'�l����cW�!��1)������ @�o�F)OC��Z�:85\|iǆ?���R����-�_�>z�s�љ�������~Lj�uKF'� �,\b� C�K��q�ZY��V�/^G���n]��S�s��Γ,i��v&�Iq��������粦j)�S��k\��7x�����%���R�/�SI�H�iB7o���u�I9�F���N�>G����Y���u<e��uZ	qh��sbˌLG�wWՑ�Tv�#8kC
���]�R� �w�V���9�Z1G���A��?2j�˻\���0
�|qК{k��� o�����v���??&;�,��,7jz_��b�`x]:��5��e�,����� �����A&�q<:v���[ɀ�#��9��H/�<x֙2.�M*g\���T�A�J�+���Y�74\L�XG���M��lX�>m��r7��* ��������d�*��OZ�����JY���CYS#����ŵ���!G�d�f\P�+��P>���B��8�a�g��j�ڎx��4G3�|�I��P�JЌ�\�d5�x���Z���/\K��ᨌ}o��]����	 L�N�T���sj#�k��y��fM�w̞)�]E14�v��
�}{��̋�Y�C�aw�L�9Iu�G�N����g|^��J�	�c�呟��Zgh�f�\����k�,�̅J(b�?t�O�'A��̇�B/J�]�z�ςF�>0�����H�nm���_�i��2϶)!�V)� �e��`�P�zm�b�w�7�G���࿓(����gf��U���k)ex�؋��mgS'���nFElv�f^��s�Y,m�&�8����cb �?g��Z�CAA�IS�>�t� ���ak!ب��MD����X9�Y��}��r��DmG�e��B4x�X�8E�C�v�P/��M*I�X��l󩢬�-l>�+v��Hp�.,گ�=OTUܢ�n�^d�\6$����^�']!�t��*>Fߏ������R�nژJ��_�V�.��F�uBǝ���黃&�N����
<{Lx�x^ooW6;H+��5c��%WO[_.���8���e����*��O��>bL�տ��z-��F���( �s,vN� e^��㝭N����X6Hxi���]d,�F� C��M�����	U(�<'��Qg|o���DS>nh���lTϹU�'<����� ǖ�m�Yp�Z���~��.���3��v���`���8���C���E�f�g�j�r������?�CZ�`���}c�\n�-3{�*g��lnjâF�J�Z��q�#�d<&`S =��#�4$ܷAy�N�P�ڮ@ [���d��8YE�*��*G�4�Ezb��I{�S�AFP��M�Nsw��ÿ���¨��z���Hv��9��C�O��?�:�o�g
x��'P ��A#������:�����i�v@",�l�C,'0�d�y���� ۟�3��9� 5���+k�:�YYU����6��u'd���gݳ".s��*k����H6����z�,�<b�WrY9�����n᯵�?T^+���#�ǄtB}�Ƕu΄�^�t)���|m���P���;��	��Av@��CR�;�������2(8[�x؃&[�	��FD%6*�k3<R����!����)����?3:̐1a@Q�����XyN͎U!`OK� њcZ�� ��(��"}�(�\PQ��
0W�)�Q���y��*�i�Ԑ���r�@�!u�`"VS�»�+�D�����T���Tl��i�(��{�v��������R��T���&[	/��Fz�ߨ(0K>�X�Ѵ���Y?�3���U��S�߫��
&��]b$���Ow��a֡v�!~����i�����6�"�����f���SaOĕ���&�9rH�j-(�a�}���^fE�ux-�xQ��]uz�e&�ʡ��Z�z ���щ.��'�.�$f[�u�*�@�3�t��ު��R��V�.U�ʐ{%��yͅ$������x2HD�d��V�6�����H�uN
 TW�˴n�0hA��!\�F�7��J2��6���P��'�-˚3ok���#>$p��%#*���ϖ|��~D��^t����5 ��O�
���&�0������!�Ɏ@�Z'2�Eؽ�t&�j��.��waL��ݑ�72��n��w5Z&{9/}~{��F�A��L"Y�.|�'6��D p$�F���\��s������=��
� >��\jH���F���З�㈝��b95^�ǉt8�>[��Õ��]�������*���I��YO�~������^�-G�vM�Ӥ��:����i4�0w���}fz(���mdڠy}�;U��ݵIȉ����d�8�$����пG�,��3BWC�Et����?X �����0'ĕ.�t�
J�2R��Be�+H�j�<>�$ �q�f^�^I0�pn-��8]�$�?��9}B��3���ڻ��[�`���U����2������QT%g|ܷR��A���̺.�¥Y�i:�6������V���O̖�t:�t-$�Oi�6���#9����*��8]�ږh'�ʞv�m=h�j�[N8]V�����6���T+��2�q�9O5�@+�`O��(��}�B�����ݩ���B�M�b���Ę��)k�{Vv�޻�*���F��6O�h,\.}�k�����q0��5dg*Ǆ�?��^Ë��� G���"�*�O=0J�i�h�=kz�t
�H56���uU���t������݇���-��
̊�ӟ(l����]������]Ȱ዆^�m��q�����	�N���9�^�n��q=B�#Ec����-���vEO{���䧴���p����z���7,M�)��0Aܣ��=�L��3ݘXL�(\�#��,L���H�L��j|Q����6=���>�_<8[��������_J7NK�0�XjE�<�ӂ�T��	�BR.=+�ڳ�6zf?$1R�s���NNGa�<��PE*F��¢-�6�〘�/���}d���|e~6ѷ��F�K���bH컠���YEO���������"�����?�0aB�����{���Κ�bv�G��y5��xh�ݝ00DIs_�Q���y�b�� T��ҧK��M@��;%b�1LG����U�=O�Tͱ#���#��N6���_-jVM��x��W(����o�tj�c���4K.'W�C!@�NG#8܍�.�]ε-
�MT�FX�]�X�O���p(�3寇_V�=��R��BX�V���9նO��#��Xdb"lvm7T��F���c�R�T�TE��l�F���C.L���!#T0!��7��}o�Ic4:/s&mt��l�����L7�u��ެboE��:"�އ7 Ff8��u8@��jM�T�9GD�Ҹs�}Q�t1<OB�<�6j���ȊY�M��]��w1q�'qP�����a��v���!��zu)`�8 ݻ�,gJ�Tg��p:�H�o��w$���x��5���/Mψ�coIN�𗓇�>x�`fJ���帊��A�aLl�S��8i� ����8��xl�71_@W,�,���3��6�*����b�7�L`�� @�����D�~����#�i���Y�� �kJ�S�H1Uaq����W�0�y9��V /c�yHj�G�b�-.ޡ���0#�G����Q��]��Je8�g �+�yc�{�"�\�p�,Lж+�=�}�Eڻ�j�$m�Fc���]�����mYXX8� ��0o�-q#k��9�&���G~H9:N����s���<�dD���@ݏ>�v�~����*��$4����r���I[ۧ�-���P3K���pM`�t�������)H/�槕��i����AP��9Kg�)_����Yp8R4dz\�m���8�@�=toy�8e�Wq��K/Ւ��m��.B:�+�Ȓ7?_T��h ����P����5@�v$)���1g	���������9�XV)`���P׉�Hޢ�s���⭢��t+�Ӳ����2��3P�:�$�BF�|	cZ��(C�cjGR.E�R��N�T�K�ݿ��k�<��hh�&��S��6��d	r�/�	͌����a�%L�Ȋ�So�����o6�l����M�R�h]F,������˰^��<�+K�Q`�f����jŮ�k'&G�2��������S-����%8�ؕ��?��j
nJ��R��R�ޡI�e�"���8��N�g༯����%&�n���ҙ���K���k2�B^��n���X��,z{��ªg���I�tEd�};Rp����	��;=�^�C�)��B$����V�4(x[[���ð;wm�P"؃b囥��8zN��B�n�	��QDan`�F�浥3�*����J��]Pٟ�*j9�ό =H�	�T:�f�l�W��[AN�@;ٿ��s-��s������lW� ��4s�� ����u�T1l�pu&%��9_9Q�%�n��)[����������&�2�NZ�^��k\X���ߵx*zhXQ0�{neW*�#A�	�����M�)߅ISNnk��z��XIÒ?��u��*'>d�9�p&B�g��\��F�{��ؾ�� rHs]�ۜ��Z���h���f���'�]�N�zh���k��Hݕ���o@[-K�{z�4<G^��7������ǟ���
���/N)�Yp�����G_%��E�J����fH4��S"^�� }!/�O�Y���/:�E���.�궢��f�zߺ�*nCZt$ �� ���x,�hܬ�Nq3�>+ű}G~i����H[������F��ا��f�^�\�Ӷ��W\nc2%P����S*�^M{��Q�F._�%}�ć����U�6�O!��8$��8�۴V����]��j��Q.4�����&��E0�#���R�	�\�����.�c����֣�d��igTu�����S��Y��	��Z`@�w��{���$����	  �/��qO"͊�G��6.�	ĕ���B���u��:CsD�������'���2��Jbd�[�݆�ǅV��T��.��Fy(�~�?'�z84"�Aę������k㮦@
��Q�a��>,�06���~1���o��tmK�P�t:�M��qsr���k1L^D��~��Yݠx'��T���惥����y`r���4�]�r-��vϱ�r�f��6�C4�t�[MF��\��#�n㈶��L��
�o��,�>y���zP:Qh�1���)ݑ�>&��X��|D;�u�����\`2{o#�Z��M��U	���'��`��Y��W��&�'�ݵDu����-��t���~G��l����fG݋�}/q�>N�� �*�缴)1�[��N	Hh+ )��a 7�W�D�/��lj^C�a��M]��b�m��P܂}�MTf�ɻ�wJ��P�i@�1r�;	�2���nr�|1~w����h�����,X8�������k&N�8,���乨�_���~�X��H��Z����:h?���g�N,4�sv��1u�C�37YmX7J��J�4(9�e��/��)`�SC��ggM74�ĸO�61e4�;��,~�PT��K�^|�Lr|c�~���x��C�Y�h��-\�fM��?���<�B�P�'����,d��r�f�Yz+IU��g蠝�ʮ���m@��dI,��7��)`B}�,����p�c
# ������AĿ�|�8���.��I;���eKl4 `x�&$>��7�лS���6�p�j�!���3���mi�����|�"�h����1>�	�M\��hf��[I\���.�`k!s��$�yd]"�D|��] {<K�e���)77{U��5Y����'Z��2�ʢw��.��Z����3� ��v�۫��_�<���^�d��f*,��9!��WJ{�ݎ�<Dg��2:�TiD�Nj�'�L��,d0�L�R��þ���?�����z]��9��;C�*�b�]��L�	wl�Dݞ�A�w:�����l`	t�*���K������9����H2f��{7C�L�Q�y��שx��\�Z�}\\�\_��D'$��#��T/���������An~���G�L)e&��QD�6�c8���cfO�j��2��Td[��<O�aj��7�nIq����57�B#x�Dqӡ���eF��MT�^ӣQT��1"�Ŵ�\�6���p�"P�Y�\��F��KVVC�:$p�;�;�c�s�\��י貄Ԑ��=.%?���FO��~����
8|q�;��R�pd�|Qm{�W��9L�ǿ�������F���SN�.�p�|΢G����)#�8(\K g��JR��3j�* "N��`���멌�4^�.T�h�[?m�*�i��q� c�&O,��vb0����/��	\�n�5���֜w"�I�
��;U�RgU9z=}:e�!�
Y�e��	�7䵩����z��#`����Ek�)թZe�*3�mj�-�_��У��l!P�f#5�b2*���XSy��:�Ê�!�t03CB�d�T��EW�I>N?��ЎM�vY+�Z^#� "U�8������c�z$Gd�U!���hʛ�ϥD)gr�ߣe\綳�g7��VG���$������1�2�R���N�
��.R�����إ� �Ŝ��d���y�;���$�y{�z�$��,��2�u�K|;�l�0�w ��4�r�
�����^WK?�?2�����&C��ԝ�pQ�t�̄}���sL�_�[��'r��/��ly�ts}}7ិ�\����A'}�u1��{�Z�%rW�z��k{93vL"�aB�9gkc��	���A��B��ʬ�#���{�l����J-�-c-J�VĽ�)�>���H,)��'���͜ĿF��mb�5�X�YV����x��Q�ַ�v��f�+��O��!��q./��z�^�N���c�T}��B�F2�Oy�#���q)u9����n�1�$�Ro+Ϳ9�z�ju��l�U�jBs�����G���[�e	h�%�V�N�K���e��=�D�VHGݾA���%�����Z/���7�+��T�!"����I��9��M�}%�wpm%M��O��Х�h��5�U`a^��٢z�!B*� �IA	���,���U�C�����)�~ɣ���ݶ�˜.l&�i/u�H��/���3o�<.������@Ϲ-�N�R�?W�-3J��!Jq�lյ�:�tw	���,^z������������$:��5��~�Q��s0�H����=��ܝ>�:�US�N��g7����!5J�D��2�+<�\DR,�~�r��t����d6�T~�.M,��m��))��j  �ƴ��p�4�y�<�BPa0�*Hs���7k�<�J�%��XƄ�i��z��(�/5��Y�c`�18�ɻ��j#f�~D@��p붅�>vu��Ѿ|��R���!Kh�c}88��R�`а~��P��[
�"%�?��S��Eγ��]Z4�i��>�:p�AE��G�ݥB��B���`�矸ǽN���w��#j�tXW0`�V� ~�yg�Abj���ŔRD�;N��dM	~�$z7c%�2��C�w��:���'ω�u�V#���C�C<d��<����<��"w�/�b0F�SnA�5����/T���5};CR����a���}d���OF�!�����L?����� eْ�k����6�K.aBO��4�:��͈:��>G�|s�¸kC��Ì({'�ʔB]U_U��$X�8Ӆ��]� �t�⵲��-Z
�� Ȗ��A:ߑg;c��cjᵉ�Z��xhoE�WH��t��t�?�.Y�K����>dC���d�>���))�5}
::���/U�3챀X���-үz�v*�#Ii�~����F�7�<<w�Դ����@�X>�X�spy#"�{�P���z��ĉy�gӆWx{��[.!����~��Y}�^�Q��|����8��g+K�@�R��� [�t=C����<fjp0c�D�g�ԃF�,�U���X���v5r5�k�:�dı�|�:�����;���;�B��'�7�a<�������>ٺ��o^�J(��ӫ����#�&����(���v)�ɛN�������=�XӰF(�ָJ`^ba�S4:㓎��?��mg�=��;9QdQ�ф����|̸���
*%�?�0� �g"��x-#m1�~�>F0Jbjf������J)Y	�����7_�i⽵�p^Y��Ϣ��0�Ac�t����BxK�����u��I�ć�W���V%t�b�g�Y3����TB>�s������˦�߻�u��s.E���0FZ]�@����dA�t����6��G0!ڦD<�L�4f���
RsT�(��R\~�vJu�rĜ5�K0��{�l��|�;�k�Xf�q�ٿ�[ߢ(�=�ҬAk�?���`7��x@p��<���bX0y�L���P��x����[_p��&���ʏKs�e������8y��s�X����iݸ�ځ~�l�on$P��-�H��:��S@����龄#������S���'A@�yDyj�����'�!:	܇��4��:+*٫��.b�g���u^��ƪ�t7\E�B�@�^�<*��H}E��;��~� /~D��VD�:g��Gl�X�AQ]z*vE62�Q��]�	mD�x�o	2�6(�;�YHX�؂�n��MɜBF�I�����~;/����'g1�7�Z�{�ԂI3�b�O)w��3��H��7 h-��.���gP��_�y��H#��jy~E�1�4��g_)�����@�60�������ŉ*�bY��m�0��[ X����M~n���g�J�����1
Y�.01rdY������hڀ[IP�
�x;���d�����{[&��6]8)Y�w�V��
:�h
p�xCX�*�ǌP�Q�}��(��u�eWYOɓ?"��R��v�Rn�L8�K���g����|���ǉ��8;���IiD��V9,���5'����?����8��:@;iԤ��B��+�.���J��~$���!�Y;/uV�܎Z\ȃ+�7(u>�q�w���䫀�����o�'�R���y�P-��L5D���ߟ�B;�ݾ���9��Հ�X�MB�qMP��.������M�#�v\S�4�m:hO�ꝭk�?���2y��!��[ƨ�L\�� �
�3=�=bI�T��g�͔���u�̐�̟�2BmP�*	�Jm�Hx����x��s���\�)�"h/�0���X�VT�`��� ��H)%H���c�0()Q�Wz#�	v;up�,T6�4�<hS�%(cF��h�cL�u������a!M`�b�$�r��'љ!"�eG,�������8-�O��&���b���A�T'+|��
R��6u$�;PW��[>k�W�yh.S�n�z�_���V�Y���ŭ���`�9�bC�̘+3  M���	��,e��$^�&��v�p����	Sb�sh���g�.
.���@o��oJېE�����4�ɦ`�X��L+Ѐ�'�;��Ǡ<���lΟ�\�U���e��7'�ǖ�<�˽��|Ygo ,�m%�?+�.�<ր{�$C�02��c?�WқӇ��t�L
a])X̻�V4E��ػ���n�Ŗ��{��rɂc7�>�f��`�&���gB�@����ZZ4��
	����ụ�ɪg�M��y||g�h��c/�4��t��?�6㳾�Dw��:!�j�w��u�{�Ͽm���TaW��b�9���la�ֲ���:�I?�
����Č,�A�[�%�;5a�"��0�Sg��n��q�������������NdJ�ڜ����y��Y�pOz;)�%�V
Vp����ۂ��he�箣-p�-�p�;�&1���\�$��
]R'�[�T/��6�������+t
W��w#r�^bkTvB������� f}+���^48BHHU��j�ZZm�u�(�J޼m+W*/p�垴�Kn1:;�$}�WŘ��ݾE9�C�p���J0}ɉ����ȱ�޹t.S��T����� �?S;����zP�������^����SprH(��z"�0�,9J��ؤ�=��h��U��s�[Jn�ݭ���!�{����-l�Q��d� �9���/!r��k�z��j��I�<1��cf��E���n��0����4,���ؤL�i�]�I/��Xt[�G%~�W]%1f2"��sZT�J&���J�q�����a#�_�0��#��z��K�1kW�Ӭ�@�d�J��.M&���+���'▫+�W��Op8�W��1�K��zY���O��$��'���%C���0%9���h&������)�zh$�ĉ����I��6�e��	�Gj�|o1V�`p�&(C���`�t¥�}��Z��t�蘪
=~��
<�D#v�?�dN.��QUL��VؽJ�p䌶jE��
�Y�Wet�چ}	�o�,��\��MQV�?���[ZsW�UAU['���u�1��9L��s��i���n{Ad���ߘ��:b,���������R�4.���� K�`z���S�$x�l�Cr9Q16�J)mؿ�xcտ� �����i퉗~�x�&\)����[�ԝ��&�TO-����{<A����sGa����N���e�N��o�қ��m/��o��Huh5�~�agq�T�ܤAe�m�@n1�1���u�y��m�X�\A6��RI�5�7���Je�p��\��x�*RT7x���g2�5����C˵�M�/VD�ς��zVe�-��(^B�����Q�45&U�)���xx���5SA?���2X�8��at=_!A�[&W���61���|��>-1����!�
��瞿noX^���(�
�h�GŧkL&cQBc&��ҝx���*)��ho�Fg!��%>rfz�4���������j�q����;�h�vY/w����b/ �2�竈'��ܐ����O�-M�K�������ʰ����h���E���H�o�ة�{>��i���Z}�Xyի�]әh��Ww��H�z�!�aL4�����.*]UR�]�ZR�6����?�lxf���� �Mf8�8 �L}l������Mz��5�_Ս���OH�1�j��#�1�����#����-y�*Ȟ���p��	�^�������	#QtfO'GY	n��MJ��$RS��8�B���`�̍��C����'%���P��{���c�wÈ���Ĥ/�)�=+�F2�<�1�z��op{�#�S3�#�3�÷�l�Z�g�(j�wS������G`��v�p���$H��ggc�����P�=?���&�Y�,Ȋ��5*��eݿ+=�UyO�Z�6��8�D�Ԝq?I�R�I����G�	n�������:�;ԌyKf0�&���;�l ����ɞ������*�������"U����i�#4|��l�r���-����v^
����и6@4"P��*D%|�R �z�'��"ӋuV���nx�+�ꠥ������y�	� �.f�1�V�_����H�#u�@T���-� ��t�u�F��1>i�ؖW%,"I�����}�������QP�9*��g�ʓ�z��8�Kw!�A�B:ZH��J�7�x\X�	�'c�v�$_�׭T��#�]�E� �%U�$Ke�y'G<�;GQ~hՇ���M��1��l�+q����M�=��1�~�'a�f$V��Q`m�_���I^])�Q��՗�nG����Ͼ��]�㭞~�4��[]K�v|Q(���/pWG��� g{}��_e��I�e-��U����l��[��>x����Sg�g�Hd���e:�`�Ƭ�F�!WD����h������>j��;����]MF�`�6tiw��p(�B��b*[<�D_�JlcB�/�0i�E��bڷv:9-������oL��D�7��9#E�Adk��_v�@���R?c\�O�cPo�c���h��n����j1Xz��!��:R�Rɹ5���w �PLm��n<Fg���U
}2 _c�<O�o��;�𙤳�i�o�B���[�!��'"�&�v����/�UN��D����ç[�i)&�	ۆۣ����AqJ�6-���R'�FM��F2-S��]�>���>D�þ#���Z.>΋]�͋�۟���|	�x��ŷ¶
UOu�`2�L*,�[��√����βB[0$$�V0v�h���W�2�b��p 5?�tg�v{�b�:��7ɒFಔ����"�2;
��X�T�r��M���P4�����!K2V�<P���b!��KwZ��}��Kj�h1�3eT����l$In�����_�Ґ���6�@� ���`�gɉ1�x�	`���٪|��acT�=��U����A��|*Ui<����&I���h�<��/����N�~�����O)���F�5n)�[�ѥ:}����7�u�* h��+*��f��
��}k�H*�c�c��G�+B�g:� ZKs ?N�5�%����\�ɩ�ў0t�\6H��J��w����Q�!��E��Q��F���ʓ�B��tO;�!�5u2LGN�I�q�a^Ex��t���R�#�4z�G4���`A;���o���{���ۿ��coY�X��ݿ��=k�y�6�_��$&���ߴ�L��Fak�ecZ!]� :*�9"#E�;JP!�ոK5�s��N I�V�2�7~�[�ڂ�~IU���b���ϟ��>�mޮt�W�A�A7�lq������i	%�zHI��~��dյ���jJ؏��,�>�2
"��mVA2h>�����/��	EV�w-�&I���Z	�r$8g'-�a9��yf�[��԰�;�����|)��2H���N�[�+��GF��B,
-��[�Mtc5
)�y\�R���Er*�%���Y�FG�1S'K?�I㼌Y�;�ɵA���I�XF	)�c����V���Z�GX�x�ͅ0������"�$���5�[xB��.�l���菠�K�ގ������{�GyJ�X�F礰|�0½�y�	�J��_܄OF�����ד����s��wb�k�_ӄ�M�{R�&��0�j1�7�.:����g(���-pB�u���G>'�ƽJ�#��M�-�W^��}ӹ�	����jq�cz�EK���Z���ahߏk�9��=�(�X��.)�#&�y�F?���ù�Bܙ�A$�ws���;Q���5�Tb�zd��!C���-�L�,��dM��^o��ćD�̊#� C9���]�#�u0�oƥy���雊5L���Q�Tc�=sX�d�*��yQtv��~�e&XY�3J����#�D�������k
��4��M�t1�Mr1��z�_x�)�g^I�&	~|���Q�~�m��ʶ�Zr~�X��9zZu�(}L�����Q�=�(Cg܀Ќ8��2Q.�������@ǥ�o�^�]�B��ɫ۷ӑ���:6ƃT�.Q�0�P�;��$Y�1I���wz���eӴe�BS����($�*�Y@�����o`ں\A�/+���([�*�ܨ��}��	yҡv'���k�)��ØE�,�bX
тQ)�� *����d&���f�WQat}���[����>��Z�ό�7�`�p���p��$�F�a &GTa�D���J����>��'�U�� =���ޯyw�_�er��7-J|� v�,�Nx�.��6G�ޘ��|��b:���)�������w���6�{t�ʌ�BY���|���PK΋�ۑ��L"�ڹ
�ȵ��-q~�{X��S�r���S�����=9�0uf?�!�i��H ǩ��vʚ�L�]���#�j;ή{�P���� u*�T�m��N�c��z��UrC�t�!K�Vo��5yfz7.���D��'c�|<d�8r�݆�n���Aʹ�<�A¢��~���o)����`2ye5ߗ�\�B�s��h�dS�Z�C���a����A[��Uwܕ��?㱤��\?!`@C�_��S���2v�b4+B���W�ot��ǎ��lq2D�h�0�u4��J�!Piy�u3�0LpE���?�ө��N�|)�p�;M�y�@�]�jt4B��O?۾߭�o[�T_.}� ߣ��X��i�W��l��h��%��U���m��e|�r�o�6ܲ�6�X���9� �:�K�o3�<���b�86����>��bH�B�h&���#���rI�W�~��O@��rLhqhz�zρ�F�}}Y�Ȭ���x�K���n{�!و9y���Z���t�WךH�N�c̌�<�P�ǳ� ��\u�:u�t�4�a^�3G�)I����v�����uܺ�H�+A"YB�ޯ(��~�>'�(Z���i?�ϱ9�����gFT���s&p�:��x�77C�o�;.�$�)�Tt�cд��jM�)����� �kI㊪�
]j ��)C��M�;(c^ֹ6%��]xw�{V����E�c�A7@
	�	��C��3ޠ�$wԃ0Ʒ$���K�?�/%�d|6x�w%ֶ8�j�i��X���!��@�Hi(��}h�6v��w��n������)zUt�z�O�����M{���w7Ўe�k`��K�@��>����%���7Y�����e�=�?G�^�?3w��ߴ%K<t�*�{�rte�B���Q��3���[u��G�<MI���Ήڣ����"��e�o�����+75RI�2*I��0�m6�H9�p�l�=C3���ތ����x�L��z�Ң�tA ��"պ�W݃��"���B,r!�4铏0y
U������GA�R��&�
�Y/�S�fϓez_�9��	T�U@����� s@�^=�
�֛�L����>��F�_t^}�쪒�J޶DT�*�T�C���Ԃ���Ml��dV�	$��l�l��(�t������ځd����Xp$[�����x�t��.~(c�0���Xe�5}�lk\��<'Ff5`n�h+w:0���s܀��^j��D����:Qi�%�
2���魱����l�������s���[y��j޻>� �
�����E������N4�Ͼma�sz�EQ[�4l8��K������(g�j����,'�N����\����"*!�*WO�f.sۏ��M<�H]�a�?g���%�|�zv�������]�_�fh��P�e ���R��?6��5��i�#�*m��'�MޖR�(4������g���N�yR�kCP�v�x��0a*$#��x���Z�r��j-{��0�䯑v�ss����|�3���% ��/:wʫ�{�%qp6%w4����b��tʗ��&�/�K��|Y��Xb��d��5�٘���Oxw��;g:
��	��Ns�z������h6���,BrmH��6}�PS1(�%�Q������rk݆��F�k����������a�k��-N$޹��t�÷��ĺ`Q�=�J˺�E�k��(f�-0�a`sq���\�L����Q%��O����ݵ{��~%��5D�p�J��C���wrzd�r�����-w��-nq�*�ɛ���)Łt��Ԡ%7�����Z�Z���@���PP6-Njs+-&��1�;(��~L�VK�'��=�6�.����g:�.cB�r��+4�V�p.����"p��M�������g^�Td�M����F���'�^x[����cϺy�� s��%���Y�EB��7��Y�Ƃ'OE�Eϑ�ͳ�'"݋��b�acZ�`~!^{$F��CR�f�5��4��4�]���j~'|fP�~�tT����I�"l�k o{���
�'B�Q��Z����?��%���O}�@��Qf���@p��e���P�hk���jI�T�h� U�;Z� ��8Ѳ����s���3۹-"Ͱ~�)]�Q�3of�b	5|8��N�lE/��/J�DX^��ЪqPZ�������`U�"%������~�ISp���U��Be>�i;��E�H��秄��;<LȎE/I�nA�O��=����bpH���O;�Px@���Z.�`&��ϑɑ^$!���~�H^r+6t% ����H�cnCnoLH���):}I}���b)\�D�{br���}d1����+��.I�2X�|�,�M��I�HЂ𫏣��e\��ǰ޿��t߰���� ��d�;@���_�g/ߣ�^�s
O�7S�����PF �vt�:���✾yن���a�N�4&�y�	G�N)���
���(=�[7ts3�pQ8�z�QCb{*mm�C�ə��(˜Չ����
g�7, !.C`���O�C���4TLZ���n/�l����0�Sƙ��3>�����D+wb��s�(��T�������36�OPqw�8���8���|riFJ��BIa�?:KQ�V"��������i��>�y�����r�9��ꬎ�Q4�R�ۗ���8��$�вy�X�T^��6��|��h N	�I��jӭ��Σ�:_���N>ow $4�@dhJ����g�n�A��奪�<��E���u��� �k�c[[BLgz��UEQu`^�j�ӐZRRx�e�=�C�>q�(���ܶ��yQ�TUgk��1�,������j���Q�w�5>�{u��d�;jª�Q��j�$�'#�a��JU�����G.ⱜX�>�@@�N�ʸ�)e��*��XZ���!`A�)�j�IMQF�p-F�3��Tq�������a�F%�O�ܟ��+_p�f�X d��:�t�d��=�2�¸�I#Ӛ���@��ܹ���]ɩ�>���_�7�<��H �z��˅\9�����eKC��%2~����b�Dd��`�j]9�0���p�;�~y�����ɑ��rI.u�E�Iٓ\ ^��)j_��%�I���њ�[�,��7[�u�6�Fa������`�� �������;��l�*~�Mھ��]���9��U�1e."{�Tѭ�0p�c�T,��$z�jn���DD�A�w�)�8�������	�30 P����	�@�p�/]�)87Qޅgm��K������W���	�O����B#��+�����p�w/
0Q�tb<`-���l@��(di�n��ש�q�@����8`qp`,e��X�>��IJ��clxT�M�s}P����gA����b:<c�L�4IůF�B��gL��O��5wz��Q"J���R�olG����|�9�hh�`���5(��h.n��W���&�m9	�/u�	�!�x�f��i?�E\�'N�ed�Ԝ�|�[��Ǌ������[����We�Hb�7Zה�_��1Aޖ�׉�[����h�Gd�I��0 ����7�:�G�m��\.�&c�;��MZ�l�@��@H�%�rH�kf��a�N�[�7�k��l �'+/�C�Y!��V�nx�JEU(�)`K���<�
�' O4�yH+���9����������A�8�pK%FP�>�� �ϦUU���S(� ���
s�od�>��8��"��C^;�I���U��~QZ-��j#�f�;�/m��˂ё0��]*�Db~�O��)/�؊ �TD���E*���̈́���X��n��3w����M[W����[s�H�� 'L����A��&~
ٱDT|��HKٯ|���G��^oZ�@�,V�:˯�lr�������m��FƼ� �:�w��x欈�C�`h�z�d��H/A�N�1bL�-;I]�c�I�`�y��_��w̰�Pzh'O<�:¹`K0�Gn߁89(D)5�7�v��R��h,yl�Q��"�ǠY���g-���7#}�=�*!�*	��<^H|��g��]�N��r �_��s��⋄�Թ�"8Xy�w �܊Kn+#{�"k�������t ���'��h;����*�I�2Œ��c�u�`�s��>�7C��d�}l����É�7��"���h�)��#G:��Ȉ�n̑�Ѻ����d�����3���Uq=ΐF��t�A���,�By���jgC���8 ��`�ߟFbԇ�QVPN�B�F)�Ks&���v�,�@��l��+�3�䈺გ:q_pzL��*�%�)�B�����wղ�}R��G�� �Rnb%-}֪]��$`��$�ώ�X�C�8�E��I��-���P��'˿#Ci7ˆ"F+��%����{6<���Hz����3u�w�j��"���m�.LV6s��/K.�Ζ�3"��E�k@k�Yx��u����	�/�/��v�$O[�ڥL���:�Y�.`ZXY�^�f�f\��}1�(�!����]$�/x�蝬{��pB�5�OhR?�J�qS;q�lm�/��Fv�_��9n��k����7{��@Kg;櫵A��$��-� <*r*�H?3�>:'��+���>0������1�̘��8��]gh�O�����U"ƺ��m�rLR8�C-��HF�P'1/@�v	WRV0��R�-��&;�'��L�i�;
^t���ɴ%���A� �ų��4d��X�{ �.�Y*m�?�n�b��g��LY���rf�i +�6�6�~�otp��J�АWS�&�:gyY��Z5�>�QDw�	�+��
c�v4�3��_Q>'�$�)��C��`5u��u��Ӂ��y�4J���iD��[/?���͹��v|�N
D"���s2 ��r�G�,�� J����&�v�aL7�W�m�"�Y�П��)X�������U��_6#Vj�B�:�8��d�T�����v�/��F��1�hq��k�Bn=�Pr�t4��cǤ��D;�jN����AM )�n��Ku�n�"�K�ǔ�՚T[�D\���>����%a~�#�;�E'?>��3/uJOw5��z}Ԭs6�#��%����xd0%��,~�X6�ϱEͧ�b����{�Q�5�KSe?�"�4/�6h�0�?�mj���Mǃet⯏���`RLq������Y�Ex�/Z�6G�'��n$�m3*�B��2+�`1|N).���'2g��Z��їB�=h���=�{}7�����L\T }�P��2ۡ�%ŋ�,�AhG��E�l�Uma����F����ԡX��W��-�gH5���y��CB�셫v�T�$V�f/�V�5���'�i|���S�Щ�:C�p�v�r���}l��^���v��H]�V85{?���2�x�,N�,�f�.��%u�oh�^&'z{�R��x�o����>q Ht�Ĝm+JQG��t�wi��g�=���.`8�q�U���M$p�>K��{u��LSܫ��������E�K��|�����K<9W	/0R��.����#Rv���ĳJd��d�u\���9>�����Rn����w����Zm����Қ\'7�����N�����꼋��ّ�w� ��#����X1�Ҍ�roQ��Q57F,�J?-wF�B ���7�9'zz���Vj�P�7�4�E�y��.,�e��b�-���c}?���&�=���¶�M����{͹��Ւ�V����/�:5}Th��$v���C��m_y��Z��M�oA+�%�M4�Q;��~��0���yN�0Ț�TY����?�ق(?�u�����
+_2�5ŏqa������O$L�cEkպ�y.q
U\�k�m?b�D�ͼ����Ϝ;7f�Uz��/��de�=Z�2ǚ���u��,� �ab�X	��jڡ/3�lyo����8�q�X�)`]b1��h��xρ�7�x7;��Ie�pC�e|��l�?�ê�� �j��
=E���#F2�U�Q9?F/Q��|w��c��0ɴ�
����E�!�Mb`r��;kN��lǕ��o��ܡۤ�r�/���{��,�$=��~���f�0NOV�s���z��l&�S��l�K5�s_��X�='��'k�ݔ�(���9��/6U!���k�Vhd��686W3�������JX?"]W���m�0Kx�]�U�8l.P��;a���RK@-	�Y�>EոCG��!��:�#?< U+����=���;Ő��FU��Sڌ@O8�8z�T}�羲.D��	�--���*��:��.����n����z��tKr�a�4�fs^�76�L:q�U@�)�F��/<(�hS�L���_ �@��w��q��7�W?������J�G���.��C�;�\�j���y��3��;������I���_�m0������:)��ݙ��G�����48qk�╧�y��P��O$���v�!�i���d�2��r��e��/9�����p8�3 ���!�����f�LX�y������r-b�Q;�ǳk�/��M�����
;W�4�c<Sp�Qp��DjF}U�e��)~������6�v�,��0�,��b����Ďh=��о���!7��'ب��n�U� ���о�ԙ��;1s�b1�hA�<恁�^ѻُG��~N�$�%�.(E��<��y�2�/�*�(��^j�)�,w_��T���q�m�QnD�X�-[8��h��uS��2 /�ՔY�ig(�7w��iJ���G�KV�4���z���z?�X�v
�Q�ɼ��t��_�#����V|e�'�CrU���y��4)���stK�'�?f*۶y��ǍJ���`��?zz<�t�1W6D!HE�5<����X�}j�:�]Z�l�q<<���b�y�x���f�־��6s�w,_jĕ��	0�R�b��W?ilq�9�g-)��+N1�1>=�x[cK����vpS��|e%*3P3/�<n���f��)	�.Ώ��Shg�8�8�AH�S).�J�FF�|3F�^f���P%�ۓp��p2eG6�C�ö8��Q<&�W�@ks�ςv�(���W�R!����6�Ac��7Mf��!e�_����+2��"7n���!�x�G[��JOV�P�N������f1�r�3h�IH�P��Y9E�;�K�����xt+��o4/�U:�/�
����x1N;!�K�m�SO�^Џ�A ʶ���|^��o%� [��>�� �r�]ࡓ�N���*��.�T�T/��5rlwU֬����po?�V-Na��4�,,s��g�|w&�~f��nk�j���Z�8��R���)OS�*P�W���	�C�����
����kL�$Nwv�z�����@��{ #W�2}lJ�Qb�G���pw��������L�Q����� �����4I�R]�P��Vf�Q-E�{SZ0թO��G�A��ݿ�.��#G�QX�u�rJ�m��,`��k�H�0�;�޸4M[����q�q���OU��	wه����؝.�B��Z��o��MIHW��?�Û��;ۘG=�Yx���+B�]5�X���� 0e�үa�uO��GbH��d)7pc)��`�F��� D˝ }�}�e���c1@N5Y�{y��9�16ա3��L�"f�B]���>��v��tbCT�B�z�R�}�����ې�DH)
�"6w�s\}û. k;��9�S��AI%�N?�y}�5k�4؄yAZ�R��!��%N�$��ֶ���Koߟ�}��k�A�v�#q$���Sq;�o��A��� *`H���w�|o�^�ZI�O�<̗��� \J%���N��AY!Sr�u6�L���@k��Q�H=�v���.H��6P9�v��	@�~&_����_`*�������B�r�2ϭ�*�>�����\�<�n��p*g�x�1�;F�RRy�����0ޤ�u��L���Ve��+ b�f	q%R.��X�.��&Z�.7r�c����M���,�cw=~��p��	�HJ  ���C	�`�9پ�6�mw#F5���C� �i�Ֆ�ʞ��Xs����#RH���ν��^�e��j26�/.&>���k�������_��ͧ�Je�ac=-��Jn2ki�w�C��
a����,F9�|i>�N,9M����j���
�?��6)�}��@~�A�bx��7	�	����o%��X�ch#K���l1��y�i���ѳL��ii����ОWn���͌�+��./�2��������^=�#ɠgR�7��x�;Sڔ�a�R۳���?���4�B�
���ʞ9��������z���G�]U�v��p*���)K!v���Iu��1��c$�8�\�^6�4R&��9t}��tK�.gҌ���d�ɥ�{I�X�wp1�Ϣ��;����I��<M�7 +��fL��x�SmN����a��E��h�e���~�v�/� z̓���Fk��TCv�79�ȿ'(��ri_�+I""J���� ����(Y�Y4 ,�k���1xِR{ggܢ�\�*��(ٕ�~�#��G���~-ܐ�������W���\�#��3M��?a?��Z+���EO�,j���&1Ogiɨ/��+D�C�Z ��E�7�\݊Ahԗ}`��'����ޒ�ʾ���h�� ��M�x�(CK�N��0��VHmiAZ^�|g��Cf�\NCd�i����/x�yA��]mb�,��w��>��Z
��IS������+�	���q��v_��ϕ�@�Y�����~�Fx︪�*F�)���4U/TI��]v96�����x�|�W#6߻m?>L���AɊf2�,�3)�>��CA�|�x�~��ѕ���:�0Y$�h4^����(��V5�r��~[�����(z���Л��]�}���{��Y5;O:�����6i������#f=w>�C�-:D⎡ ��Syz�l~B�����A�� aj�>e�ᔞ �b'��Lb[|
9w��}>U��Y	���ex�u;�U��V&U(�I"�� �)�ۢ�=@}G"�	k�P�
��vl���u��zX�11�\\�=UE>�j�*��7�+�}qjrx2�Ǧ�41�UEE%�l!��' Z�*����Rf��pge�I%���:W*�հ�B@��S�F +��n�Ԭ0�[�&��3�GFw��=�;��K�4wC�V%W�^ٚ��z/C�?4�Cb��+v2��$���ne�L�;�i�s�.k9O"Y�h튖��(p�ĥ[��o�ݲ��%́��˂�w����{���/���PSVm
�;-)���#t3m�R�iuU=iT�,�-����iPZ����D���]W�0v{�47kF�C����8-Al�0��#��9��oS���ԩ����2r�j3N�S��I�4��
7�S�
��|t_j���د��7h߳K����r�VHt����I.�f���`kQ�/��{1i���)��U:�{C���4�����W��)9��+�PSRĥ����B���C$b�L����g�������:�$�-alj��)f�:!e0+p�?1�dJ� :��u}���7���U����y�r#��{�NT'[7�Ǌc�4k�/�>/��Ԍ�����۞M@�J�;��񇈴�\Ԡ(&F��O.�����g�-cA�]2FNC�H�D���۱@�.7��s;��ޥU��ҡ�~�
�p(�pz���E�UP�>^50����A�yBیI"E_��Z�I7�Y#�|���2�/��z��Ҫ�yV �Q@Q�p0�\�|��������p`Wh�U�"BJ� WЮ�p�2ej ����C�����͐��e��D|c�$[�I��5�a��)t���e,�`/���e�w�����l�N�<3���ٛx��a|������t��2�����ا5��<1ʗ�P� F9:U
4�y;�А��Zz+	�uH�,�M��b��,�Zw��pxt��g}J��X�Y������MP%�(�*GE�0�p���o	���IdC�
zٌ�0Q�i��:M���X���_�c��B�BI�t+�¼}��a��Xp��^+aZEd�o5X�h�:��%�O����a����"JX�x+w��.6�Ǔl>A�P�r~��*=?(;��Ǚ���c����ޮ+�`�~�AV�k��Oػ9�앳��w��nK%��5L�w>��U��]�Eh��0��AS^y��x	��[��z?�x��7�j�������sP��u-��7[�����~l�d{Z��b��q�,m���3z�
��U�j&�t�#L�6rN�>���go\L2��9�!2�Q����������9�P}��>,70�*.��]��
�R�[&~J:9 ��D~F΍�O&������tw|f�w�g3`�Y\\���
4o�YrֶR{OK�J"�����Ǡn�=���MK�s����Y�9XO_hه]�XK*��0NRb���}�&�U��C{�%� �����	��L���1�����4Luwt5��0TM�x�(�;)�q��L��H뷅�?u�T��Ƒ(z�
�I���9#m��@ǩ*��n���1|Q���ƽ�ê&����-l�{�K�d�
���O��k��������$�@k��!�
c�E:�i�Ȋ��E�fr�{�f0^�i��e�}-��%����p۬���os���Bq~!�!~�jh���]C;#(vJ0`����霁m�w6g���V�yi@1�f�A����]�I\�*M�ԓ���`�B�2|o(�j��$n��I���'����Cb���L��9�L��</���C����t\����0����h���vh��r��n�쫕�,i�T��,J	�Q�0���uq���`���I�+u��l|n�T�,��A���]<B\N�*Ќ�}������Ef�rO�s�,�*�,w�*Z@a��~h3>?���Zӻ=��	-|Q�#,��٨c��t���_�|[+�I�ش�Rl�ֹ,?�'$O߻�(�"��B�H�d���K6L�� 8|�~M���8�eI�7�Z�\�x��C�o���7aX&������5$8u�UF����>؆=�w���
mz������̯��x'l�C8-
�O�_/
�;K���l٩�:�;^)p6!x`j[Zw�KT���q�%�p����ڏ�_ �O�D�!lr��'=����ow�$>��=����0!��ͪ�9���å�������٭�d;�Z+@>(�l�9@�y����(on��͞&���_�l��(��'��|����]B�d.�����>����w�N}�۫T�8I�^��ш�¢��q�)`:�,ݨ9��{;�!a���W�La#�0mKa��f$x�3g)�gir-{<��F�<�0,�YnO!��{�Pց���F�/�T����0IH�o�E�8��v����zN�j��o��4K�7��6�[R�:�v�b��Y��ܚ֦�-=>�֣>�8���K	_M/�=³��k"<��M��K<o�4]5�)V�,�d�Ds��ҝ����ȔF_ {\o�㒳�����7����P�8DI(��M��C}W����S,�4�Zs�T��n���������\[��>�́)fų>R��︱8�B�h������CB;�p��R�Z�ެǲ����a O ^��_��t����U=�]=w�
Ú�Yq�J�P8��
j��~� P���l�f�������*���K��0gUC�pO[�Z�,��ei�8^x�����xy��N=:�X��M~�-��z?�w%�2�hֱi����S��ŋ5L�h�٢�H��cK?����`� ��}�)���MQl7A�j���+���x���+MEf��o<��l(3L�� s�%Ҍq��"j݋��vR��h��σ�� �<� ��N��"8xǼj�Yl;��Kp��%�\.˘Dik������gL��XTa�����b�t�V��nȕ�e"�)��V��i�7�PjH>ZGf��C1��pC'l�������H?]/�1M?����`M��VPay}��\ᱫx��UFA�N=�eN1-�&t�'N5�Kr�.fG��W�,�S����������C@W�o���I����M�kgb�Ȧ�����PD5X~����!�ĭ���fj�ZI���eW���m׋;��Z��������� �Qj��k�#���<��bD�q9�Q����P��e�n���=�����(�n��lg����(�~���v���D�@`�i�]^�m~���3%���#x������Ať��2���ju;Y&m�w
��|����?zA
V3Y �bm��ھ��T͓�SAHm�y�/B���f^��6K���`����
6����R�D�H�J�M�]'c�d~�Gx�[sZ�����^<�8{�_�F8�l�h��u  GDi�V���lq⾢;p��+~�`\f����ރ����D�u38Ѝ�@�L�{��>�[1��]�ͱ�H1��x�M���F;8�-������f�+�Ymد�'�����	�2�@@ƽ>]#�L�WNY��d0h��
ma���d��]zJ�a\I���~\6�[��#��8�\St5!��v�7�F��O�y'���]%�i��{�0Z�>޳'eq����n�$��0�I���7�xӃ��U R�@,QН��K%I����{�U�/dG,gN���9�G��Ƥ�54Ɲ�|r`ٵ�i}l:O�%�Y��������D鱼x7I�&��g�p��r2z�d!{����Q�����k�+ڧ����9�ia�e�WvJ"�&����@T�1Z&��	7��Ҥ`�r�}�V[���a��&6iZX����P���	+���n�W�E)�� *����7+O��ƭ,-�i�z�j�<�=��ݞ�)Ϣ��z!�p�/��y�0��^9��=��/$����8���ʾ=@�S� q��8�+�X& G��T�pP��#}�`�,�H�aPh�b�ʢ+B��բ��^�AX�8p��-�	�}�5���Fxf�a�fh���Wp#��צ�����0TE�e�xbi��[����Mi�9��4�E�T�P�,S�5���W��N�er\B#�)���B����.��%���o���"N��ͤ��8����	#|ǏL����hpm�W���僧��8O�4����1�V���~�|9��\<���2#{�RQ���U�ѐm�����%�6�����4%%D/���MN��(D�<Q�X����w���,�بA����Z����ߓ���cI�Z>72�m��@���=.���S�N��qvR;Q�9��Td�G�S:ڵ�v`��J�����Y	F��Bl��� ��.Z,I���1���*�B&Ta��،�!;a�h�X�v��1���b0J
g�%9}���Z���ұ�߼}���d#X��F{���.DR�V1�Im|��v�y�ޑ�#ͷ�-%_�]�J�B=��1f�0U�"s�>;��F&���*���x���:�3���	������+�t�"�p��i)��q�����B��;�>@�t�Xp���Q[S0.�c��^<�&XB�$g"��x�4����uD`˪r��;C�4�s�p8ɟ ��l��FĖ����:\im�PV��O%z���]l�	E�Ї�핎�`�+d:&/^�'C���c�5{�!�_N�OĢb�,��Zf;�A�fxt3[��@�U#�Ҫ.*�JW���JLzp�=4� � �/��!��Q���X�nƶ��Ӯ4�����e4j��4�@�a\{2�w����
�@n]2�i���/�� @��~bH�"(�eMmq7k�y�[���,1�F��z�LإͬXSU.��*Kb�cP	�Ifo�� n��gŀ.�6�Cb�tVv7 ��j����5��q6b��Ԧ$��.yVv��q�#S����eC�;Rɴ�j��:�i����ݰ���F7���M-s�%, ՜]-�󨧧�|н���|"���f4|�W�l��K]yPdR�1�ߐ9+\�N�9P2-
�j�(��L��j�eah��ĭi{�X�pn]���T����\@�=�n�}��߂dY�ˁ��Iم��R7�ǎ3&�a(��x��I�H��MM�:������ўv	� ٦)�t��5�c�P Gܡ(8�+yE���Ȝ��'�ghd>�֘����NM���ej���Xc��wR]6�[�g��/�.� ��`�l�L��@��@Õ.9����N}���uIۀ��P԰ �o?=!Ɲi�6�w�I{��K>˟�0]�nV/M���"1�?Q���c�m��Ś�^h�f#���|�z&߬���}}fڝum��1�yѯMps�<�W����V@�2����rJ/��,����1�_dUvP�K�Ӝ)n��m�A7�y9Ve�X�_�V�ה �x^Z�]�4������L��ϝ�D��r�G�	B��3�1��Dڍ�Q���_Q�����*򕚥ګ+#��#�h����^3d{�n�۸����c(2)�
����b����'ڜ������|*�8���l�m��O.vy���d:�VX(�ɍ]�u.��խ�x^e;�,�ĄQ��T{��1���ҏ�5��@�QΔ���P�!�3����jep��IƔ��f�!��Q����ߴ�,jnŐ�L��b��%�3�E��4I��	x�s�ԛ���/g��ݲ>�7���{��L�J���9�`��I6"Pn�Xv�")�J�!}�Zj 	�hM�����M�sacuy�8�WGi�~|4:��侬�g�թ�{�Ӊ�1�'l�]�2����f̦u_���L�(������EM�/!�� �z�Ѳm�r�ݴ�0h���P/�ܵP�Q�kS+�Ub.�?�N���ڢཥI�L�|\��;�g�{C~�Q �0��	˂��޼P4�Sm��2b��V��F!r�����r������$i����/�x8�w ���H�!���t�_��Q�����~��VYa8��m�I�s�+Ǥ��L=�gn���T��mP���Z�9?ڂ��:�6~ر	NSG�RLh=���U*,�5�%)�ܥ����T���A�(�k��5P=<�+gn��e?������d�C��GZ:b��o��|�Aw���g����	*�s�°� 7����1��ԋY�j'		tv�7�.�*��dtb�9�A��ڰ�.�u�'��K�(<Fi�@2��r'(����ʘk�g��1��B�K~�Э��ZPZ>�'���x�K>�K~��В��$_B�̙�#v����d���PU���#~!rvS^$\�Fj�μ��X���I�tϞC��� A&���Y[^�]��^w��8A�k
�.F�|*UQ*�'�v�?�r��]'��bzё������j�+����P�U��/��#�(�!�iS�P��U~�[V�B��D"�p?�]�fl�ĺm�!AN��I��T��gb���޶HT�]pp�y��&�� <�W�I$~�,4��;�%�h�(+>�u�d-6��J/���s�;�C�6�&h����@s��J5�����ۈc�)o�/!O0Z����`��/�v�z�>3Mb]ܮHP	k����m�":�6���A:����rV�9&J�짥_S$-u�.8�p7L����Y(��xi�?	yh�����a�
d0��qF�Q��v��LB=V[�w?I3�l���hg�H��lv����qF���=����t�WDʀ'�1s�.&�٦oA! W��&"5U[���ZRT��Y�#�*���/b
x���H�]�L8�^�#������U	�A��p��W%v�����o���)/+�ӈ�L=�ʣқ����i$���ҺL���j����f{\+��SO�	1p+��83|:a���X-c*�8�7��Q���x8������~� \��Z�Z��>;ŕ��-�T���Lr�t�%��|l֕??5�fR���
�	()2c��1T��g�{JB.���E��Y�ޝ`ˉOup[#��+��o�j�|�g=y��"��w��zd��e>�i��J�_�V�S!(�1~�쇨���k��Ra���膝�b	�4��q;��g���L[.S�U��>=��>a���zJ��zWX����[6���%��s�Ӗ�q=�Ɵ	x��#���+X_>�4�a��}�r��rL���.'����N�S8k��q,�������К�P�2B��@�l�w�D��	q�����P��e�e�B��75���D��k��p��L�m ���#`Ob�ւ2��'崅�.ѷ��Q�6=�r��C���f,��=��>m�E��Rq�� �ߝ�ɤYM�BhR�͆ׄ���1�|��.�ݚ���1�-�a��qc�+�䁔������/�kāUHWw�vCr!"�,8w����0�j�H��,\�&�{�5$��ݺ;�{�]��S�y%�KJp�����)�� |�ߴ�,�l��&�9�UkĮEڀ%R ���a���j˙Ya҄z�eA�o�Of�r���e$/��<�m�8;@M��n�.\�
��<=R����>Qf����nL`	O�\ �,;��P��Y���=���?����4�Ar�����n��ʲ
%A���,Ǉ�/���Y�:Y4pt�2#�@�8@��Y���S3 X���S�2G,yУf��5��#�O^��j_���ŋ�f�O��B��˩J�� �`	_�¶d��X��Fq��\+|<]�u^��������K���X^�2[�#C�&f	���o�m�Ap��'���R�'-$�;C�����ɫ��r8D9�&�%�`h�v{Ll��ԅ�>@�<�]dV�g���Ҫ��`�����?��bɬ� 3���m���?�]�c����9aQ�&os�u��a5�l)��E,��Ʒ>�����,ח��e�e;�8���ט��uR�?ߺN�2��$��s�8؍$�s��N�y�z �(��%�r��$r�r�Tx�,�f9m�,D�=�b�^��a��$1�o� �|���.�.̒I.-�
)_��2��֩I�4����v���sA���{��z��k�l��rf����	�UN��q-G<Gɬ3K�]�Aޝ���9�ܝ��!c�I�;�bd>��R/���f�3\�كVѭ�u�Ӽ&�����󢥟`��J���P)zq�B;�/@2�%�A=4$�c�r��ثA�]x e�U�g����]l��D�c�1Ӱ$��f�& �B�'�h��R]W��ʤUu�϶Ex��K��qNM���w1�B�2���zYPoX�������W�9,�N1�u�G3��rR��b#P�5����s����`�2pM��R������Qe�,��mL�H��b-nV5�ɿ�Vu���ġ�m3g���޵[�j�n�Qw�_�^�%9w�L��D�������`I�
����V���s�������<_�݁���0��x���A\���P7y�L��7�D�[�Гɳ�#�S��p+�j6�W��&���+���Q�ŕ�v%�N�j��7ZO�w���@k�Wí1h��H���9��H��f2}I�U"
�ٱAVY>Re��$H��s�\�.�d!����r���<&�s��M�T�_���.y��}kq{4������`�湅���2��sf��|<��DҢ�� Ihj)L(���ʬb�:�"�߸w�E�����Z}�؋�4�)A(
�O(����Q�?��Y�]M�?Q��I3�������q+T, ���P�?U����$n�t:δ�+^���뛧���i��{��S`���|cW���I(4ފ��C�۳���:�g&��+��Yd/�����^���&�*��cƂpjѦD��+�暷��ٚ�w	ӝf�c����h�=:2`L_��Li��T���1��0zp\��˷�#�mn[�-�!�1�jmX,WB,3>��9�ON	�Qi-`�㕖�O������M�_�0~�n�&\��l�����y�ݿ���8E����A�rWѬ1��r�b"����@Q��mRC#B���ҹ�ƥzt��Yb��><~��ɿt�E��*�z�C-l[8ew��(j� �@�(�U��*G��'�O� Iީ���r>��S����k��i�B��H8hs��"�߂A��d��<ot�!9��u�{�:�w�g����<d�<���*봌��������8��t�6sT�����J�L�������q�瑦�0�jv�'�4Du�uRe���5�y��3=��b_��~v,��o���%L7����s�Gy�R�����L��_d\&t? A���+?�|=Nq���M�A��nI���L��{�__X�mI�J�S�*FW����nj�e~,Zl�;��	�M��eEK1vT��K*��֬�*�Q� 71��S�~=����5=Gk�	�K�ۭɚ�b�o��~��>@��*.�N���|��cg�4�Y�����V�ݑ�$����Ҫ�م��Cxw�7���	����1Ѻ�QLYuc}��:�[zƮs���LP-�B3��!���hŞ�@�l�"����}����W�6�]H��D������U0��k�å�?uh�W���&���-C�~�8���h?>/#W��#�|r���rMhQt�cLp_&Ә�N�E��Wt��.�@�v��qR�����h�m�s|Ǒ7��]���6�rE�e�Ky��[:ϟ�|�؜f�Ȁ�-��P@���o��0m>�� @�B�\rg~��ȸ�v_y�%��7Z��T@���h�:�^��a�}e£4v��bZ�i�p��Ք�)~�VN��%���&C��@��	�
���� ��-��wC���J�؉�3���r.��T1H^s���&C4K�R��Ld��V�>V;���ѥ�f�V��X1�?80��utOx=�<�fA,�E I�������b=�_%�CKBY��	>��p�12y3N+�m��?��	Y`�H�?�~���ņ��D�N���wOp֦��K`Sh��h0?!~�]Ш�G���En�e��L�������B"(����J?�Jj=%k��X4D����z�ov�V%��)��s!�X��+�]�!�w���r&Ɗg_@��PMd��]LV��g0̂����S����^�G�TU��;Q���U`�"���!�/��Z*���sR{�&g��6��,Mq���[�P&�H&�O�u�Z���(�zW#.vhk�z&�}
�Cֹ���YQ˜��`�/��hv;��	����j%x�������j��@���� �6Lү��=��11.F��������r��6��r�C��N?e1�Ng�0���1	k���`L0������R�aaZu��mb�=��)pR���ei�c��$���z�iL�6��Z�@G��b�)7���o�U��Nz�Z��C����p��<]%�r2���=C&c2}W��S 9Q(�X�,_=�|��Մ�v%ڵF�ǌ�8��w=vÝc��@��{Qr/��G�����rD��,�7����U=b�[�r���w:Q1�%ښ��ݒ��ek΃`c:�?Q1ϻ�.`pt��l��C#Y3��Ȝt��5���mS �� "c�x(��ٚέL�:�4p�V��.k\�g��x�����-�I�B[���ʛ?��6���:`�p����� ��E�R(SɁۂg��9�3z��'�霋#���N�G��yl�̝�궇|Z�x��'Jx��Yʉ%t�b���Ch�J�ڬT���&U�2��uI�e%c,I�𑠊Y�[�'kΫ,[�:�>T�`V�aV�S�a�����e�vh���(P�= ��bTz}G�P�f!�F�^���.�2ͨrO� X'"�_�m��l���2�oP�� hF�(|ߗ�k����(�3��-��qp��6Ϳ���N�ը�0H�.d}:ʨھ�ܵ#�`���mLز_��b��KGq�r����v%�����6a�7�[�8b�CM��nl	��C2A��mI���B�t�\�;�4�8��/�|���z��?P�G��-�؟W��GP�ק23P��7	F��)��u����$��\E�������C�`�/#���N����aK*߁b��7z�t�=`�?����y����p������m�u��`և��ɖ��v���|�,U	4d<C�ίp�7y�FqTg1Ov��� <!&�CnH1r��Db,����˺�[�����7񄈐���g�*I�4ر������|��g�[~e�ӿӛ��	���H{���d���E;���ǞNp�U�>FG�o�BV�W5��KG��Uy�o�+P�T̸e[�ǭr���2h��
]�<_��o���AI���'E�ёG��`i�6��سQ,G^6k��ep����d����9��}! �� �&:.[2!�0�u�/|o�R�M��qwQ:۬�@�]̵sP�V�An͡ߊ��;�����L�\7f�8��\z�븣2Z��K���l0d�p�������y��%%�!������e�#�d*�7�aT���q�s��6V����e�>��q�n�E����Z�mL�INư8UT
W~e�O������\���_��|Y;T	H�ϓ��8Wb�1gД7���٧�)ˣ���0�,�Hn�{�m]��a�/�1)�2�Þ
J�Jp���n��L��ܜ�2�tLK"	���Nh���D6��T�	�lD�g2�5A�b�(�UƢ\O#�N9�𼎇"u�r�X0��V9��6�����, Ν�Z����GX�г���&���U6�`l���H<?�
�Ʉ
��@�j����Ԛ���Z�A��WJi��nן�y]�e�� ��R�w�rep�ϿZյT~.��	W��Nn�w�3;Gjx�Jnv� �A�Zgh��~�D�¨���'YH���G��L�:���F���-$��m�c� �]K߿�=��~��y��&-��ѹ��CtXl�o��;]Լ��h$�毳��+<���Om���{����w�:lSt��?oT�5�F��ۅV�r�b �� l�gk���T�k�V�����s_к��"���>��|I�E��9��X����!�1�߹�-�����4�8T�cߚ�64��̭A�r�1�&��g���DkC5���י?�h�4����|�0r�ڨ���s��<i~���) ��s�lP�O	�?���?(� ����t[���5F3Ȼ�b��&`T-��h�l

�����zr%�e3H����B"z���\z7��9�q_BQ����6ͶY*��_���C���H��5rv�9��s�B�=��Jq_[��+<6!�3����/}0�W�ԌG�G>U�v�1�0~�Q!�1v�,*U���}7b�Hp���Nbe~~�n�>�7�O��2�ڹL��<ż�wՀ���9��S7c�8RE�#;����t/��cƍ~%_���C�)�`�BQ�U��C��P%��1������
!�����>�YX}�4��B��(m�l�*�0$|��g�io���a_��\��'ؑ�bG��<t�)�i��`
�*��X��L۸$ID���q��l��T�;�"4~�p�z��}���'�,�jGM�򀔧8Wt�&R-�.�C���׵.��+W6��-Cjy��I':T^o�(/c�S��&]bNxj���.��=���l��+�wpO:�c�@Ă���KIzN~�Qt�#�
�|:���m��{�����J������>�׿��GV�练�Z2P��M�2gۦ=^8n}P(ә�9O�E�viI��n#6ze� ��i�eʸ����e�|N_�UtXF�>+���{Rj�/X�X+��|�o=-1�r�����B�݅�]�8(%�`K~��;H��r2�g="t@�u�r5�75�����j{r�X
VS��y�hH�e�>���m,��Y�Z]������&4�*F~U�_��g˒?���G��U��T��k�Ц���j��u{O�2��˯%{yh�!{���~�{sjF��T(�`v�& ���s��͆�c>���6WU웹��� {�{���I����ݦ����
!�(��ã��Ԑ�&��x�R��vGs��9�"����j1z!D, �8sZ����^�T�˵��������|#,���o\(��3cЗL�0�-�DT1�j�D������س!�}�z��yM�YP�n<>��"Y��U�� ��$f�b� $zm��-����N�[���.�֢�Ib��93j�B] ��SIU+����؛F�}�xy���Mt!J�u�_���0N'8sv�A�"��)��p�w�������w�|w[u�>zV-�`�k�4�5�����q��/�^�HV{�}�����J�� �p�{��?�>'g �-̨�W����$3�2z_����
�<d�0��r�@�~����v�+nP���<6=5��H���#=�L�'�E?���H�^r��֮j�D�փ!t;�^��ӆ���"���nep��gd/�O��/&��
��);7��Ϙ"7��5�ћl˕C�bxc�(��X�3V��c���),C���lv�5 �>Fq3�;��>��m��Q�mZ����#��&�R��G��&����v�yGa��iB�W��5f��U�)5���%��k��r�Q�>���UwQk�X����B�CW�ɔ4f� �i���u��%Į�d|�ӯ�K�H��+���o��3���}�F��-q(��YC�5��g���:��^��Ǡ����^�*)�O�8P�+�θ:���X��)V�=����B�R� ����:��)B�+�L9���;A���t�zla�k<(��.d��H���"���W;5��dCG��~��86�X1�8d�W*��� �}^��T�`7	}d��˺D��xf4�����2:���P�s���������)�3ȿ�,P����l��}v"�$ʾ��l��B�h�+WF]�i�Å�A�ŝ}�O��%�\�Y%�P��2�Z����q��h���<F�jb�!����[�z��$	��+�����߹�j"h'��Rv��=�WQ)����%8^)�!� �A��k1<B�7`\1;����������b�ɅM�`� ;;ǨC�֞G2d9Fi�RL-|����;80'0�@����A���n�pS�
7���vG�]�L���P��6p'*�'U��Dۇ����CrF�U�p,JV(Zr`=����G��DQ���ĭ �_���JVx��E��	�%� O�w5@�NX���rP^
rB��_U:����~{��:��ڠ�-RY���v6ڞ{�T�q6��?�2�v�2�����\>���c]�پ���!Cj.���Z�O��s>Wb�;�q�я����=}����.�������A�$R>)����\���ML�	���t��B<������
��F[caǭ�1І���������I���`��5���J�@��#o��#�T &��q���8:���'8�Ӑ-,��W7�l��s�	V�-o��!up�L�i�`�,A�ra�gǨ�����nt��rĚ�2��e&�-qt��V�_$�����"���-��q"r�#�G2�sĂ�c�-�4�|� �2���L��=:�V�����57ZmÄYX��i�́Y��Q�;����E̲Y��#����`@jAt��Y6�Ӫ��'������v{R]�^#�펁�Q3�C��Ϩ�⨘��R���w9]32��7Z �e��JOs��sD�����x���+�[�$+���'��E���r[ʿ�u��8�����~�R�����|U� I�Ψq��]�����I�W�i8]���j��Z��+eLh	y|���M����r>�<��l��e��K�T�pu���翯^b�\v�I���X��xb9J�	O8s�ҁ`xß�OX;л.Vb�든��)fl`���:�6YIf�°?�k����n�׌��'dJmq�;E�JeX���S��u�j焄k�B	i����H ���D�P�R�1�:�9n�E4�����|"cs�[Rh-H[�➻Q�}���-�|N����}n�@�v��E�`�k�� ��*�7��qı��w[2a{%���Mx��mrʺ}�8xu�w�Z6�	�S���D���0�S�?�M����0}l�;���h?P�Z�SmiI%�X%��%�h4�(�y�V�����-k��3�VB����D�E��f	��@���u���6 ����������D���z�HJ�r�te$;���OJ^���&b%�VQ�hYkqF5CC�ZB�a�8�6C8�K9o�$19��g�k����FjK�����Eo<sl,p2��7i�o������T�4�i�Qj��s�dԖE}�R�.�ky`���C�@x�v|��?�
8:� ��WB��_2{��˭�G������t��{��^x�!� ބWwiK�Z�l{s�ަ�= �ߟv
1k.WBzi��Nȁ��QXfPfL�����'U,����+������&Qx���$JW{r��k���X�%�-O����Xuʰ~u���&7��j���i��ɚoe�r!�w�H!J/3�b�S���
�rnr_���N���]	9�c'$��)�e=P�Z��#c���	an(-�r7��n}n��
��b!S��-P0�N�y��dz�;p֬��M�A�u8��1G�|�Lc.~Y��M��eã�y`\��O�-�Wl�~Iz5���s����jW�I<����Б̜x�PC8�d&��}�P69�S(cOY�s�'/�>��!����.Nm䮍*��Q����������e\���{���_���ɒ�'f���x����n'�VMe���H�� �m���ӗﲓz�r��2�������^2y�R0�6���`׫&4m����� ��X��m�Ժ�ʠ�,fP�)�P�=8.�WG�/Y�2���C�E��B���F�f3$Tqn�;��v��1�:��O�3m� ��죓��o+<�V����C��,���e��I�yg� F�xIT���>����Kц���8`����T6û��%����hI��Ftυm���w&�EV�������&hJB�䮨�5g!瓼��X�bq���@���W�"��'��sU�L޳b���� F�{�ë�N6������襂�'�����]}�����U4!��S4�z9�K�I4�}�$��1��s�y�oю����\�I�6���L`�l�"{���B��9XH`��7�Q���S�&(F��=K��IB{��O��p"�N�!T?�6L(�D�c�$�_����_�h�biC��q���bE�m��gX���#'�.���H˿J��L��Lg�T�oX��
�|d`��>f��
9<	k��)]��BK��h*3}���O�xc1-fC��xj���!6I|\=���)��l�_����%�S�b'�@��]yQ���\m��Rh�}���ђ=�"�����;�����t���LeK�v�O��Z��+����&�V��X�~�hZ�p��a����G,~�m��� �qK�ƞa��Z!B=9�1j�ka�M��s@�b���S)[5�
����:��.����}��z�M�/`���J6ïU2oQ��W�:�'�LF�U������4J�j�s������I�u�N�?��,����ݫ����}Ɓ�.��ʗ0k�j�?�l�6I�3Ϝ	\�E�(����1=Y�^��H�`���R��V�Də����pi$�ݨE[30<�x�3�qiAP�L�|���g�2A7����l�^ې��'Fu`����^R�L�e��a����BMF��-�V"9�������؁�,7�,�w�%	Q��&Ƿ4��yt�ߐ��A��~W�N����6�R�츅�t�OM�ȍ�""Q���H�Y��&�\#�����4Pp>%���N�Q[/)�h%`� iQh˯`t��D��ޟ��[�aY~=+��$`d���#!���֔�dN�P���|�`����#��cx��jn)
�e[qH��-n��/*��I��PV�=�o��8Rp�w�A�ə��ޟr�`Z����z�Qn��'v`���1���I\	���&�W�OC���{Xk��*h�wt�G���#e����=¶����IL��:I��Z��_�W��uuп�J$�RM�LR�����!-&�)iW#+	���b+���`�����G2�3�k@��k3�Z6���`TH(�h?Etq�mf5I�h��*'26/Qg���='�6N��g�h���W2z�i!�CF�h�ȱ��=�i��k��)�z����F(LC����"�h
G��*��� J����W<�Gd�Ȯ ��gb�}�j3��M�u�ar�Y�JU�hn02��ęW���,j�J[�M���sT� �3�d%z�l�"eB��	�o�*c�'�� [�[�"���V�����#$�.�����d6I�b�$���/��o^?����oF|��H�>�ρ*�7��8�v�D��؇'\.��c�O���]�V@p��1��2̊��"�i�ґ��̬@�j��C+E m��SC)�[��YJ
��.��:�����R~(2sę4�:�\�\����c�p�8��a?�w����Β�����.�*��q#c8s0J�?�Z��H��op(�<�	���e����c]�T��Z�;�q��@��3�.�J��[�)o�2�e�3�<9��E=��p;Gb%n����7�+��b��@Z.Qe\d(�U�(��θ/�mO�3��S�{}�
��[�B��I��8@Z�jف~	&9(m�+!�ܕ���eL-��yL�����/�W���̚�C嶂��@��H��8����PK��Q��������A��`��z��
x��ҽŞ}�R��m�w*�����ޛī�_:��r��!��O�����k��E~]D� ����W���g�VWjL9�Ե�#�/�8��:���W�r~6L4T%�=qh���ݰ�~��X�@��,8(ʭ~�jV�g1H�éܠQ��7
u�G/	�X���rgg����6�ڳ����C�����筶dI�VNV�?i�F�F�]g�fE�Cw��]�/`t�!����D�J��s�铨�r�L���Pٴ�0PqY���<;K�����!۝k�9`�B��~� �[gO6;�x�xJ�K��kJ�3��}�,"t�q)�)�,�q�-uӗL����C����rb��e(��s���pa"R�,!���!�F1Na}h��oQ�����]*�z�I��ݨ'B/�#�Z�燃��y�Gm��z�Jfp~P,����g��0pN�2Y�X�oJ�(�W�u��DJؕ�HbR��',�DӬBۈ\�^y�'�n�����/����������g-�KD�V�$�VM�UI�9��4����V�"?e�181���;����۵���y��;�uڄ�F(��BJ�P�a!O@~��h\ĵ[)V� 2&����U�$v�=�����"���jP�KH�i��n^{tT�3�����2.���F���F;����,�I��@�H�JQ!�l��d�U�Jo����a� .^��!"���$X�ry�}T@�b5��)������:<�Ӻ�M]s������]��-��eU%�@N�i���z�3A⫀���E�zj��69y�m"e=��ϻ,J�y����k� �[�}��V�T���*������T$T���Q��8�h�a��5B����`��A4y �H��Lܱ��J���G��̼[`7�H$7���e��a��چ��IBw����\ZA��}@K���۽U�>dp��)����!�u�}�N.�r�b��6@ZDHQ]CH���j7�Ι?=�G@>m�Qm���^*v
�}�T�Y��T�9�[1�1�1���2�5���Pc<>���KEK=���6��q�W6]�9�W�h}EdH))dw)���-���o�Z[j���I�-�7x�M��+Ym�Bq���Tl.�W�(J�o?F�B���SCAK!X�y8j����D�9��Of,���T��Y�c���ܝ�f��_
���x���ڞ;�� \�([!vhE1<���_�C�%2?�-��+c5�����g�vCP�4��h|f�%@��q1�t��?zBսx���	��I�����Wdbpm���X@�!�۴=���|-&���uNP����ܱ�Y[^��ޙ��]��t��a7Z�����<  8��u�q�x��k�=��&�����b��g|�H}F �'+�_{o�9��M߃x��	p�6_�
�Q؊��HކC!��< ���yC�;B���X(V��X"x���~DYɢAQ�eW.�	������ك��g&�*nD4�.ל/TJ}.�"�}
����dw�I͏�T��`����"Mi�"��X.:�(���Ј�#��2�!i�D�eY��+Lx�����J���N���f-Wĩ`щ�/��M졕g{W����ǘ���r�����p`h��k_�����uՌ�,�-e��2&� |����Z�rz���U����y	��;��s����E��9Q���ڸ��mV��^�X�O��v˥{�b4���C�TQ��cGbR�^J��lj��8��!�q9���z�ۄ��b��K�L4�� ���?�Rfg4�f�Ymy��4d��b#��7�F	!M�<i	'm.I �M6�42�Y�]���fOc��Ȭ�9x}��{����a�E6p����L�<�x�5�,}��T��&��e�>�����nFmV�(@���F�t�O5%ɲD��
�g�i�s��׀G�2�����Z�_6N$�B��C�,U:ޟ��{�m#����b��~$�	mw�Ҏp���JT3~�7�,��u�0f��bFj��-;�Y������.�)�CbQ;���}/��M���*O25�\?)�Ј;�g��?~$�iwO��64�2X�@�YB�K���7��4�^�c9���$2��2I��Y�����>RFS�rZ���'���V���Σ3|t����H�1N#aǇ$S�s1�j`��q�����1Ңy��� �-�wT�����m��x	S��˿���P��I���v�F/5��q8�W����0G]'޸���6U��̓b�\=eK��`��ԛ򎩰0��2Q�7�L�yr�-W]�;�MAJ�#E��w�B~?��&+/ ���L��;|��=�(��N�v�&��H���A6�:��F�r�?���u�Rj�6+��7��g��(q2M����1�/OG��~6Ϯ�+�f����Z��岭I�:Ϗ��#��s{i�w�����p��1�x�s[l2ŗ�T�TC���1���PD�F��r�C:���Kv^�:�C��}���{�B���� >�F�k� �֚��-^c��GW4�
�b�Z�f-C�@v%��U�.3߇�/�+[��Z�&�9�#�q�5���\�{%n)��t���Ň���@ݐ�P��5.��ڮ,E'��g˼���	s02�Y�)��ώ1��T��TG����s�g&�XL%t>?��4U%��O�3�8���]�E1Μ����rQ�锷��3y�g��8?�ѝ�'�1|
Sd�'�x�����ړn��$��6��~��?m�Q�@HY�z0�ɝּ/���q��>\��&�3��@��b_[ט�i�^Y�/�A*�i�o�?w}
�+g�Lԯ�j�g�؇[3�u�p&v-	������[��>����ⅾ�B�ku���rl�u�>�N^�>I��l�?�J�1��~:�[��1���:g�4�6ÅX��>�)�d�$T���[55��'�$�>mc�?;��XR.p'��V�T��N�>G�b�_��߾�H�T�U���J���-�}�P� �����9�$P���ӹ�/@����!��#��W��	��f`0N���T��?�zi�;�����:Ci��7�u=$pi]�U���.j�Z�� ������֫��ˊ�L����q�K_����#Y����\�[!�ϋ/~�2J�	 �Z$1fi���x�nR�o�eK���]ۇ�Y��M������s�t�I�:9�u-ӕ�GWM���i� �i٢�!�Ғ�r3�z\]�pe(�H"����&;��f�]�u��px,��]��Ux��.���2Xc�3j��"�[^p�TB��8���|�ys�zV�Z�6��|���-׭}�_5��
$[�]������gٴuY�
XO�Q��G�{��e��g"�d������Z"axiA�L�5M��eh�y��MI���
8�o��<J�!S+�I�U����݀���Z����4�����e���!!4��'�mw�5ŅU� :8�~�¥cD�����/��KZ=p��N{��o{�x+Y��V�좫~3�p�u�_|�*SE�r�!���'�S�/� �p��U��H��s#'x�6.K�52Ιt�$d����^㣙�9r������-ڻTY�l)�K�����Bn�\�E1�g]0<�����ZYK5��S+�Gĳ�Eh���3Dv�����y��,���x�R�`�����G�A@?Qӎ�����z1����8b�7=O������,�Bk27��'���k\�/�8~ݷ�P�A��|����\q%�5�2�ޔ���-�X�PQ�/X��у�ˍA3��z��	q�82V�I��S:Q�RZ(����(��q[IY�٬��{�U���$�7��П��)v���~��[���>O���A�<����F�,��a!�n��ZlJ��{�f.˯lBg���Q=��3;iY����O~w-�C�%;�Ρ�|h���o��aT����o����n�˱���g��e
±���{b��+��Y��ZQ���/�������L��t���.Ɔ���MN �
��DD��Ko+��7n�9yĳ����C���э���Ҷ�ۦ�Ǌ�(e�9*Oo[��d���'��+6�=�gfhV%>�����5�R�sw����@�3���	�8q�Mm:�D�V+�øf�"ϑ#9P2E�rheX��tVn�^�t5��X\*�g���6),�5�ܠ��;�%���׆�5�M�H�m������C�+MzW�<���`�<���*��.�i�0��N��ؘ�������4�J,��[�6��Ԭ]�j4����������I=��0�qX�ʎQ*�[x7J��I�'�TVS������Z�:F��|�x��y��<ٞ��|�!����W���f�͏��-����I*��ߔd�Y�f#�Uc,��N?��7��=�u�ܵ�ـ�^�\C��%�2+��MN��8����z�g�8O��5�0Y���=�2�wK��Y�i�L�߷.��˶T�㞚���y�N]M�f�A�����.�"�����{.�::��p��K�������`ѐ:+n���ܨ�\v���#̠�f��f�G����C��3��mG��4%�'5� �Y���%/���Bش�M���?h2� $�$l��1n,�z*R�����T�T����i-+�=CO���L+Z�zn�����C3��<�J��vD56���^�d�<53�Ē!�����ʖ�;W�ɳ�(��b������*r��o`Q�d�� V��.Ӷ��|R�Z�a��ܱ�����+E*?�{ <����@y��O�\�χdG�w�`�[�/��GI���)K^�_�R#� �4)�!�_�!�B�]�)2��t�Y�'^*t'�����.�Y��Ϛ��	27!@�zMϗ��&s-���Dz�V*Uy߅]o���#4�_��8�K��;���QNk�%�'C��	G�K�ʮ���n�g�	��� U��ߗԫJsYhpduQ΢��\�7�u�RY,<S�ŉ��������L�ʹ�Ƿ�3p����k��[�Q�k�:Q��cu�� y5�\�
�Q�����f���RS1bC��n��u��~�r�)55'�Y�GGPk��Zm�6���X�2D�! �-)�v,�.K�.�3�cm�m��l�Ű'6�Y�W���|���>V�j, n�$`�bx'ԗ�W\R�qD�~�5�]GY�o�l��_�Eo3�&�&���ӂǴ���(Tز{��R��#9�T��(��L4��Jy��wH�d���] �R�T���z� Q t�\E���z���B�Bc��-�.o�g�����1a��<�{,�|7�6���m���+����F��4"�B��7�/���^�N�,tհռ��a/��YX�D�-�hl1�Z�&�X�C�`�� N��#�D�녊���	)a��b�y~V�=�4<h0⥁>yfn�phH ���}�j8�m9V�<lxU6|
��k�p�B�uBdN����qM�$�	�)�m��Q8�+př(�+�.k������|��p�����Zs�$��t�� ��M%1
��L~��Y͍]tՠ�8#�[}j��PE4>ގ ����Q���X2��`�F��A-��yN�p]CU���&��)rh��_1��nou��͚6�Dx��ڟ�2=&��!
��*�A���� lF_�~���2	��ht��܌�l�����z��T��Q����\����Q�gw�7��q�u��a{�)|�3o�jݳ({j۳�{^1���wk�t��������O��ˎW4Rݳ�m5��k� R6&�:�����}§��o���0xc���5�O�ԾBz���8ZU���v-q��$���+�Fl���a��fLG���Z����b���jU%�S2}kH�/�6p�7f�GSڌ��|�^��&,T~}:�q`*�ԏҝ���5Q,8$P~7B��谭A8\1x��X��.Р�ݞ7Z�Ȕ\�䊚�!6#��Uٿ�M~PCrMxK/���3���X� �7��j���S,,�������(a#եR�V15�Ӻͯ�m(����D"�m�r�������@jM'v	=Ҿ5�,�������7PU�ں �f{Nu|I�p���(:$�e��%~CS�ˠi�ݠ�ˬ�;�h9S�ءL����Y�Gl ~���1�G�h�),�6��p��bV+E��O!~��prR%[E.�����d�^h����BtV�>v9�V1��lo�d
jfJw���ëѦ�(͕�y-��գ�j',�f����\v�K�*)o�A3*�R"ǝ����\�/:\���WȦQI�0��:.?Wf��CEoiQ������M4�����B離�R9�ny����L����%�k|�M�f��.=|d��\ѽ��"˓^���ep�FA��ߥ0�O�|���YW�N��$�/�� ���zG���@���B̠�qڧ6���`/@TW!��a�Lב� H<kE=$������yi���4�U�����˴q�7/�!G,/���E��U�u�TE�l~��kڄ�껒�N�����q����C�������KA���a���\�P�硚42@[�(�/o#ʠ�FO8{y��F�%�3���V��eu(���Q��%�U�d��&$���+L�1<9��� �+�m�c�Z)�1�~�֌�v]��v���C@���#gݶ�g���Я����m��Ժ��>��ҥ�+���cK�����}+U+f1�#��qJ�Ձ��R.�)��;x�,�88b�[��Q�yb6��w��į�\`� 4K�	���ݔ��&T=gG��t���]S�����\���)�Y�[��8�D�k��a@GԸU�_�K��=˟�H���O�?�dј������K���+�V�GZ�S�[��u�&�q��Zx7�l@�]��n8��}�E�p����*�� ����������u�1,C-�ְz��V��A��yk`C��;��X������{�t�?!�W�6v���Jˊ ��s��لx���Z�<4��^��k�u�:U�����ag|v�l����K `�4ׇ�/�G�:� �;r��%k�⡸t.��ۨs��R<ž@��l�E�Y�Y���g$a4|�
����U#�:��5�C�C�$�>X�M)P?S���.��Ӟ$�̬�����<����(zv�>�[?XKO����$�x� �%����M�Q��6T�Ψ�������v��p�'���ё���
��w`���}�r��E��d{pe3�U��;�A:�:HA�:�̀�ʔ�=B�ex���n��~�7�"�#�x1\�w�e:�e���V��# �����Q���v������b���EM=Q���WDk���ҲlPz!��6�3�.L��ɵ�=�G��z��mYZ���<(ڋ��t�;�����)(��n���Z���tB�mxF|83ZUGuۣ�'�i^q�Щb!�jl!���QG��q�H�Ct�.�g�ʟ��1ڀk��jB�ɑ���m�e�[,T�O����1}54>��o������N��?&˖�+�z� ��?�� �|ś+�M��B�mz
���o�����-�D[��&���(k?�Vk?�mh�g�VyU8�!,����_w����\�CS�0��5_��B���=���Q~z��p:.ؕ����Z)�v�~�q�<���m�e@���'�C�&�����h���$�l��29D&�~($��_m�=�7G�y�&����'����<qӔ .غ%�R�O�S�Rӑf����P#��r�0�j�3.���
9�Bj������slO�)��v�=H�+��o�,O�m�#Sb�F�,��'=b���iY��]8����}�;1��cE|��Z՝N�$��"��w��	.���}=JN�n�#����3�w�����jrH|���	�4�Z���'A�m������osF����XR3�7�^��P����"�޽��۲�4p��ݯ$;���W6�[�ʟ+֦&6�3��:H�2��1 ����x�ko� ^ХVX6rr����?zP�	j�A��-Z]�|xVr����[�_�v�����k�ɝ�5��5��w�H�T�Fp7�R:���� �{U�9U�2$�����n[� #���.�?��4k�E�nY?>b�����&�*�dH� _��������Ҩ"];*Lo�î��o=�P=��/$�����O�M� 3o�M{ᖄ`W��t���C�A���������9MG��\�7�d��rOG�ge�Ry������']a��{�+o�t����䈡�T����Vgިr���79�h� Y����>�����D���5Ѹ���{��7��VO4���'�,�H6�g1�YFe��Ӄa9L|c�Rji�(7�S���R�۲9�G%oj��7���;�Rke@��`��:ǰ�6�	Zah�"4s��#����g��U|g:n��KW��9ߴoO��02�/g� yt�Y`
����oX[&.h!p|�Q���
�nn[�}�"�a����Qg"lu�|K*�@ Rl�*�X۰0�{�r�ȯ������{��$�4�	U�e9)ݐ!5��$B��P���D^B��l�=Zz��x7�N�u]�Ij��p �F�)��6e�u������M@;7��1����ne*��2��qn9)�������s(J�(y}x
�Gss�]P2�8$ZyĂ
+�=���3��Q	��l�c�Sl��lO�bk�D��%o!V�U�N@+6^�����6��w�U��L�������iͫP�d�*_��ݨusz 6G����yL���qx�%����!Gjb�uJ���!��q�S���W�O�<�$��.��e�w��Z�\z�ߑ\�d/��wv���Ư�aa&j��ߏ?�݃���xv�*.�n������&��i���u���rj`�S?os0)��G��E�@��z�K~�겕n�NZ��Vu�gl74�?�_X3v�!�)�<|. %^��� ��G�r$����e���zBѨY����1`}� ї}��+�T�ɨ��94D��޻��m�2�#��\���R9�-nґ>[wN��b�U��"�I[�����1��HaW#J*�A-ֹ�xF�zxYS�{&��4b�j�2L��;^��e���֫)�9E���v�՜J!.�$���Lzx�?�W��1B o��t7;��xRp����ᬊ�b��QM<�}׌���+>?��9��F�[I�r��%�`ܥ\�����"�1��p���u&�3+�d�2�#Rej,�����)l-�����4�Pw9���1�Ib�`�Ρ�nP��WU���n?���I�������cq:|��~���V}�r����O
9�T�ۥ����5�Ǫ�Wk�S���<�ja�c��g	��C��"4�86���n��<d�iu!i��
��h5�����B���{
��Ma�T�=�3�f�0���������@d+*��1������ـ&(�r���5ZK�Kq����붦nnU�zW˶:Fd�o��0����R�N�kl�߻�,�r,�_��!���G��~A�7��1ZZH�佹d�I�(��*��ҹ��N;�'I��OG~ɓI� ��b*J x��k���4v��с�M�){%ߦ�̪P4ژ��u�݊���Uot�וG�/r���M*\���N���dDBn�M�q�ei~j��/aO�f�}�=4zز4���Ԓ�a0Z<�J���Q�K��T�):|* J��=���CX��4n٤ڿFUW��k�%�n/,f�h&�g��v��h��h�Hp�(�yoX*�f�� �Ӈ����!=~��{�* 7DG����(G��@5u3m%�%mR�'ݷ�≐��S��y�
��w��r$��.���\�Z��V-4&�C|�Z`+�T�!wq@���@̬�ΥO-��"��1�Ғ�.t�.�xܲ���F:� ����Qo�#��	��#�l�I4������=:�Ԙ!�N�z�/�gP���15�	0���&p�p��<�0�P���F7f~���vꦍt i[�-�G�������`�7�J�)���(�L�V��&&�V��Q�����$�� �QR�C:�Lu�E��]����{.�E2 ��fh�5n\!��(�N�T��Ƽ�Ժ�"���E��38:��3V�$��6v�O��B�\��_�?�4
��v�ŀ|�֞0.&"�AM�|��+ZɁ��m_E]ȓK��ER�S���N��E9�n���;��rK�}'c��O8���Y|��ӆo�k������1����;H��ư���bo���yJLH����RW�0h�W�'@e���U�f�E���+��RcfR �~4�nEwF�w����_�4��~a�{��M���{ųD��9�h�3��-��da���B�Y2���DBs�2VgΎze�FČ�4`(Ӊ [�L;� ��>+���]�YU��V��Ok��z����V[�c!Y�H�+7-b�V�;?� }�Zd�{�:���-�
zfI�t�ͅ����;����?~�{u�C���%����n���� ۛRts��0���`��r�E��.���lh�Ĳ�U?���N�U�/�.og��7���<0c�5�Ы�c�i*�j��6Gb�Y�OM�9���p��h�Gw>���q���x	;���f������a���GT�Ȏ��6�n-��p�J�`�~=���I��n�'�/�.�hA)#�*{�B;�&RP����km���@��Y>��[���&�B�Ɯ��33�.�|�����3S���]Έ�;"���;n-`l�?��@2z����Stĥ�܆�WӸ_�ѵ��2&t��Dp����X�l��{¶?O���l���ܧ���{K�#*p����W�̀�K���f\*��̍KjRރ�߸Y�`:~��y�Q���H�ӿ��fJ�9��YW���ȴ��C����'�QNvz��x#>-�|���W.�U��� ]���1?7d�V9忛�e�χd��/ƳQL��u/?f0J������P�3�H�HƗJ��y4Ƀ�=	]D+��H�N�.��&9�m�U�W�P^��ڻ��\�"[�?�$�|�΢��ftSIP�p�8?G��{-�=��35c�r�V����4��d��_��`���Z�S��x��RZ#)gS���Ax�ͺ<�/!n��3�ݑ���Eܦ�������ن-� ��6��c���W&�v�2r{�����X��#��=.����7���f�y5���9�A����kFzX��������4��_�	 ]���7�ً�0�B���sH�ە��닒lY�]�3
�ZTW���A���ky�y�Uc�àu��$N�J��is(�]q]�\#lL�w}���)�M��`"�+c�t-��x�V�z�� �v�ݶ�=�8�I��w��ŎH�����ӬjO�"�j�@����sh �^`S3��M}�,aoF1������D����C�:�(J�9����~TM!��^�4 )ӗ)�x<'��d@;�^�o��~Vd�c�(���U�<�A�b'J�>+�j߅.)8�ux��z;V(��j}�)�I5B���i��U�^St*�_ɿR��Qi���ӿg.z��3F����TG
Ԍ�%���ʼ�r��JC�G��5.v0�m1�zסt&E#�I��� ���d�"]����scQ�L��*�iҷ�^;�\�Fg�)�ZɊ"u��kqIE�`�8V�;�����(�����8?Y�c͜��d�owCNqD����τ��%���Z�����RGh��s���X��<B��v��.�q�_���d������!�m���1*-a�Gb�4���OO��]�7�]G�u���K1�JZK�r�}b+��.���O�����˧a-0�V�)�\�������=)b��wهI[q��
��)�jC4��sYY���ߓȿ�{jI��5hy����\v�P�}f�y�RjR�T��Ko��2��!�7��u���uYH5��`Mh��tK	��b����%����r$�SąoynGXx�<����������{F�I�S^���vNvsbM+9n�D�}Y��:��/��-@{�`'��x:� �`�bRrVN��ץ�� WLJp/�dH����1<�[�D/5`8� �ݬ�ߍ)�aJ�.�$��:��W��,6i鯔�C�^��Qpy��U�!\H����L��BK{���M�,�ad�N���Zq<��r@P@��,���V�xQ�}|��k�D��p��;�P��ಋw�ԭ�v��-���|���w:���
r~����0��As�z�]�čM�����Eb7�R<\_H����`-*nu[�9s����yV��q�3��:��AM��^*D8{Wr��%�>��ل� �L�Nr��자�"�[��򘻣:�>@���Ni��S:+����{b�\�.Λ,����y0auT�r�Hn��8e��H��)6cf���M9�A��.�c��E��ӵm��[��xu�2�Q�Q-�$j&��F��7?Z���,�ٝ�(�Pq���#I���.�v�M
iz  X�����@���]7��şգ�Y5�E[�-�נ���7�w	s2��e��W�>�\�_�<�M>ȃ��.��4�-���sKc�Eoޝ������a��$���۴��y`���x�����p�o>jz���th�B�AM}���У�~�����9~�/�PMM!1f6a9��E���;��j�hw@HD���Bֿ�/C@2��y�#����h�K=�i|�R���!�+`o/%RF�1.'k��_���&�����9��4'h��y�5������lݷ�G��4��+A*+�_�y��K/E4OK�}n)���%�x�@l�!�̫�;R�����:.�b�(��i�3��L��;��'���n:�K�u�'S\D�J��x���&��ɖ�N��H����3�z4ץ�Z��	���#� }��9��=?��:�l_7��$P"�I#�#H��S��%?/v�{q4�e)���p��+۝��`7��϶:��9���R����/ř#sz=@�W+���r��:?��"k{R�H�����B�~��߅����"`!Y��p<����2����A�}�����h���А&�)�	b������KЌ$��V�!�;�ҟ����%��@`�(�D7�1�5/�Ak.�ga��brzA���ۧ���>/ϡ�ҏ��R����:��G�<��=&k�j�1��$���x7��%����ę�`��?��#Q,�iP�K�a�;F�}P�q��"��/\�a_@va��O�r<�Jޗe��_�ǚ�	B������筀#,-�mQ�����\ʜlxc'|�{�r���M,������i���4T/���`+H|�7`�s�o��L:*�l>��1�B��#�s� �~ɐS�.��>�Kۘ��J����tt�'i�/W��RpQ��z���7�d�+�J�[1mZA�������خ,=���eZRO>�NŨ2��4{����N���_��h�����7��d�N>U����&��Sx��E }A�|��#���Ba��˲D���$z[I5��%ф*%hr�����F�sL[%>)�ܒ��-Wa/�k+�6�����vW�D�G�db>�:)��z��b~:<s�4'	���]�Rh��q��'ZUKN�刹�<�P���/�%^��g9lv<�-7�3KgPh��P����!ٳΧgh�Rɠ���X�>�q�9÷�1}f�� �h�k���>�@��f�H���l��G�6��T��)|��zK�hUʈ�6�)wH�%��B�[�_-;��K�E���Z����h�����:� ������Ƚ�ށJ��J<E�5�F{��1����a.��_�LR����U{��Gf[jx�t�q(,3&次ŶV�3����ՠ��(" �q
6)�w.�E3��ʄ���^@飬J�Ja5U�y�yZ&�>�n���uH����`��C�1vC�B�p������	���=��ؽ�XRU�keF�������'K�c�i��Է�/Q���x8��5�&
7&f�`(@�����_WI��Y�g�$��D�N�BlQ�4z��
�����G���)[�=���1�s�����-)O�+vŅ����S��z����˒d�Jx���IU��s������hQ`�'�%��>��E&E��U ~�F��Z����zYptU y�f���fyl�'x$
�(�;,�P���/�o�c��C{Q��b��H�z0(��hBEb�G�X�jT{�ڜ�ؾ�{�H�fJn�t%?������@*3�6��-�>`�nn�
���S�f+A)�vӿO���q\m��=~��W ���"ۉ}�ل3�`���=Xʃ,�8�K�5Y�5p�9t��޿��j<���zpNs]�����5�<X�qʲ~�ʜ��F]�j�iZ�^���ޛ�l�B�&_�Z��� W֡����R%?�����J��^䍞<���<xe�d~�r��ku%4G^u0����J'3��I�#�j���E��ᧆၑ&l�_��٣�C��=�5�7������&[�Yi�4Nw�׍?�uXP;�`�xYRP˘�DC'�&���+{�p�;W"`���y�/��K�
�Aް���/R�Rο�`����?橥�;��laS8���G�G�׳��g���	LR)�������'�������:�����R�n~V��ϕ���
��L�5K{�3L~�������ۏģ�� 2X�T�l�m�@�h�~�28*��LS��_n�3l�B;��`p�I�Z�ј�]�T
�*.�H)�Z%��s�ֲY�6�_����V���l� �q�� ��c^t��������W�"���9��D��eG��ˆ>��e�˴L�n��)��Jz��K$n�2{��t_ĭDVm���X
��l���1�l�>2
�jO�o���4�"����܍�%�`�h�k
�ۣ�����>R�?��kl#U�N�ژ�G��@x� �����T��ηү��_�/>��{q�12��H�k�� Nm�����D��a��ym`!�m�(���R���ܐu��F��ӭp�6�t6�:P����4|�U�N=�u����kҠ��Q��d����g=?���Si��]�����]y}>~t ��;��!̞^�xՒ�%�#�"�6���Y����j�� ��K��Mx�|M0r�dd�ѦXi��@/�2]�fcNz��,�g��W��,F]�����[!��D� |�ցQ�?��d��a�ER���^��'j���ݭ��᢫��74��\и��'�� ��Ւ�<�>.�� }st���(6� !����Y����1N�D�^_Δቤ��J��I��� TѨ+ڔ��nV�}r�X���#�!�[�_n5��oS	��?�����sΈz�Ƈ����d�cǽC��]A���ۅ�O�J\O���H��R���Z���tb
�:�v( _N�Ɗ�+r/.*�[Q��cTH�miؤ��^)�3���#�����{�zf��p(��m1�q�<��������}Հ�Z+��_�\Y���_�@Oa_�� �ro}�WQ�"��w���~��z���M�����n�V�@�\�{����t��(	�]�:�%�����y�Zcq=n��cQTE�Á�6��:#意ԟ|2;A[�҇�7���'7��!�����@	4'z"�~�d�Un��mOŕǪ	ydn�*w5��ͤ��Е
���� &p��,�W#_�5zhM"���i���p�:V���p��"�]dy�Ķ���`����`��TC���~����Y�1��#E�Q��Q2��=�9]DCsS�bM��O�X<�
�L���ws4_Ch�*XZ�?���{�������r{��s*I�*��B��HĘ�'�A�8�Q߱:i�W�j�ԋ�W���Jgx�H�Ԇ'�X�
�@���0�������/ /��hV�J_y�%��������1��v!D�Z�Yff������&C��*ӹ�|����2b�'nQ���4�4�|L
ޣ���u�.�o�c�_�M��]�N��)n и�-���W��З�3k0�B�˝��L2Kf��o�C���cU�:�fI�Bd�F�Z���M%�N���O8�ym�b�e�߆B\�h�T�j��cX��>F��D+>�_[n�گ�s[�*��_�7TA�*�z<\kg7��Y�CO�+�|d�
�3q��W�rR�Vd���;��%����S�G��w.v䎆��ұZ渢"L`���������!WL��^w}_S�k	U���������wEbީ�t`+�T��J�i��qX-����Hfm�w\����3��u������1Gб�ps�b���/���pq&`v������e\_D9%*QR"$S5���1|�߃(;�9]�D�����H&u~�Y<8����?��Eg(���I�kp,w��y3/�m�:�(�z�g�g����]��-����)���CxƴF;�����<�(�q�!�6���{'�3���g�����`$�7l.�<�������w��Q�7j���~��f\��4��8V�̊�N��'��Aiç��|���pl�Q'K��C��0�٘��Yh�!#�����kO����J��z�Y+��"���)�'��
�ǐ �a����f�0�R�n/����7�4�XD
�Jt�B�� �D��PZ����o'y?es�Y�	� �X���au@͆�8��Z�-����Q������W���M�~4�`F��2���/�^�G��+O�ӷ���ߓ��3�yp��g�
��|0�F��ψ@>^��l��fR%"��F�b�N��@��<O,�ʩ����vl{4W�''�7��T�|���G��Ʝ;z>ɱ�/���f� ^��=��3�ɚ�꧞3��
�h�J@V����ro�C�Hסf},ɜz:�����!���4JOhM��:���4=��ӵ�^�߷�IӅ�O��QZw;�}:������$��q@�M����vV����)Ot���[�7r�g�z}��BCRn!���4%5[���������1y �m�gP�{V�<��v�M�N��Q)��D%K6�c��S$��/p���I�=��k����|xd�z�-{I�}l���t�an��B��/���:�t�p,B�ۣ��6e��H�7��=�Pp?*V����*���,j���^��=q��F��<���N����
�Ľ��B+i��c�P���d�}�En�G�w�Gx�zg�d�M�%��9fY�ad[y�vHᢆ�K�N�׶ob��\�vU�ٗ����$��_��H��X}�VX/�l�_�$��R�j�/�h���݀�.��Th�=,vB5�r�˜�0�m�d���.WL����=�ǫۧ
fjjQ�P�#��ыϭ�2��T������h�����s"�7ï��͛�g�G�}�~r6��!K��d�@�lP��)B��\y��6bB8�(��\+-&���7�6`�{j+r���mE�A�O���^�G��d�����=�[���`��Qy��LS5� +�E��z�}z{��t���"���������S��9�i&0i�0���؛��
�7�+�GX�V�g<k�7������`v^�JIj�О���;Y��M������,ä)�q���{uL[���Fc`Su�UgF��$��w{�!��)9�Ljv�a������\p2�9}���o�&|��7�ӥ�J�Ax��@�PiB��q��6w[��UsR�����g�=�zA.6E>�,���V����y)_n�sZ�fۦi��z�B\��{�cP��ԑ�YpZ����;H��J2��9��.�1ME��Q�TL��2/��b޲�}A�T�?]_U����#5j\y"�1�i.$Ty��Gbc9p�YJ�Q�e�:Nxv[('l��ǵ.L�A�kd��-�<��T@:aM�01eX�5�[���7ߛN����̼y�����Vry�7�iѴ�:���K����C�z`���~�������A�^�Z^ԝ&��n�Z	4q0����\�B��g��`�'!�Iq4a*���qr�q{4��t��k��:�t@ED_�}q����p�#��̆�]|n�
oa��g;�4f�oz,�E?�>D�.s421).z��Z^ր~����M�& V�^s�r��������_�QRpW�|���:�=Ls����ٕZ�K{��ӱ^�����2�^�v��Mr�[����;f�PJp̓a�U�ƎH�J���f��I�N`IF�/�e��Q.$�_-�I�EZ���דjE�W%ߍ�{S�x@���P�<��v_��:�X
u'4��6�BEg�ƈy�	zVht���7׬/q�,!�]��Zo2q�Gx���@�(6,�
!~f��Į��Ir�]�ᮠ-���Q<gS����Al��D0�'Z��^�޳5}��N�e��n%:�(�k�
a8`6��o.�A}z�/��[5�>&���Lj%�,}b2�)��P{u�(��!�s~�����ርuW�f+V>x#���j��P�аcpVz��iG�=�*�&2�܌��l����'d,f�o�WJ��z������=�o��pKvG�Dq��ҵ3���o�Q.v�"{�#�+5�ImW�2�������R�tD�`�b*L�Z�tR�(Ս�P
�.EąǘWr�]�A�(�y�	`��ƈLT�M��Sa�+{�p�I���!!o����X
7%��D�]%У."ې���RN��ܨf-��cu�f��5!�AS���.B��bq��&����}�\��Wm�ߖ�r���0!���@YN�[&,_KX;}}f��Z8��g;�VH��6��IE����+���j�na2X��[�.F R�����"��W��H핒�p��G�ƕ��`���`��Ĩ2�2XY�h��9����..����g�wV
�V|�
�(&���I�[��>F�%�<3��������Y_V�)�AT�]�@Č��f?�C��|�|u�w�ص�����$.�L�l�~C�-���]���Q���k��;�^V�.���V(�j��#�0]��H.tҤ�!��xEԶ��=5xV]X�ex�R^�/��L��)��p�,��~�(�!��ԣ+ٴ�
(.��i�)y�k�z_�̅�!�7-<��դY{�kb���;�mZ.�YEy"g�e�~f�	�%�@��\����F��V���޷�N�L>*�I6��[=sր �R���bT��h��Sdе��bw��ׅ�z\Zn��y>m����9�e#dU+����i2 !���ŏ|��@��V1�ծ����,���b��N�q8�=�B��TM�S���I���!�r��C����2)nw�%��~n!#���JIj���f���+.�Hڄ��bR�PmhF��"�t S�W[��BV�]#����һ��i\d$���e93���B(���B�pf
:G
��a(/�3�Ջ��eXIl:�`AL7���_�\)�*~ux"�aގ���D[�Y��/�t�!
S,LC�3�����3�h2�c��'�Fu��)i`ts�ũ86��2+���Ǐ��}h��"j�c���g�[Pu�2`:��bq��U�����<�/�L<5M>nD%��&�P���*0:�<�FR��`�#��r���2qc�e9�����`�ΧQ�ʑ��Nt��A�)�u[wG�l��w2��g�O��4;:-h��%���s2�4�H9�%�R�*���!�'!�I�e)@y��k,Z�N�-2��}.]�u~����-+�b�Hz�6]�&��#dK�Mb�l�?9+����	��֟�9)���8n���� ��F��Ι��gX���Ǜ�Gq	���i�Xm�f��^��`+��!����0S80Z	���Ȍ�5ڀ8?8k�qCby�∓���1��OA�j�^e} �S��E��?�m@���F�e�o>F>���у�fѓ�u�4K����k*�#f��~nx߹5�V�)ff��7�;Z �*~��g�F:��K�&j�ڌ*���iO���>��a6[b�,Q���ssu���2��K®����jd0�����#��7�"�7�%Z�,���U��т��j���V6cNw�d�,D�z�:<�py��������y3�T��p��<	5ǡ�O6$��nyh̚=V�/�Δ�[A(Ω�D�N�����DkU�㐃o�3]3�W,3|:,6���V���:Y��S.)`�A�P���L���4$��X����gE��9�~yb��
v�[�f�Oc���?*Z��g���؍0��P�*��R
arκք`���1Y��ɒ� � 9���#�j�>7������i7�Q���)`��y�"���T���9�]��|\��"��SH��C.�K䔘��	�N���Gs���hH��7ǧ�+{��6
��r�����
06��8��u�?�j6=i^����"����O���j���K��w�
 u�L�����S�j̙ Λ��ߨ1��n�y��~��s���W	-�G<d���"�ޗ�w�R\�؍	�d-Q�ˣI�Z������3�����������}U� ���[H�$���C����e؄t��yV���;�ڇ�+�@��WgDH�=9Q��_�N�\�.5Ih�'���M9� x�$����  C�  O�M�E;����V�rO���mrc8�"
�.���wy��	��T9���L6c8<;�d�����+���}��aڲ�j��sj��՚_�d��8ފ�yr&�7]C�X�ӌ5�/KWi�&�'��
)���'h_H��SeR��^_0KX��A����C�?0Ư�9;fA�X�Ǜ֝��L�g;��S�`>M��م���w�H��;������j"Lv<ÿ���YlK�Z3@�??��1�_����d����?Z%�3T�ع�����Y;U���]P����p`z�.P�T�zKQ��=��1\�De���bs�>���A��Z� �$��w��$<n�i��r\���ݎ��.���p��������g�}�7��n��߅�K��z=ʮY����l����"/��Aue�NLP��8���P�-忖����S���o����Ba�C;ډ4�L��^���6��앶C�md;�߄T��S۝��V:���p�X�$b���ċ��ܝvq�͈�X�q�XVS���˯�!����^��S���!("��?�/Ⱦ����ZtLrM�KŚ�����Uj\��c ��x�D0q�,k�~p�n;���溆B��d��n�YI顥P�~0Q�%���vc~\D*�B�t5M��\�������VD�$���i`����oLd�	~�a�>|h�w�"�J��/��[�c�qP��^W3����w�p8����e�d�/&���& ��-�=�7��ǽ͓Х� Z�i�!]����d2��4�+�����@�\3�֩M��^�ș�p��B�D�ҿ���5�^���6��n�[v ����6GY�_C-@#;�Z:������GRj`{O;�A�&��*ۣ׫���0�n=�y�_��T����^t��wJ����e��)�z�rg?#���j��2��9H�W���7�k��w[��1����C�A�5+�b��pi7V��|���4��
DA����bZZs�Ҁ#=���Y^���*����y�k(��%E�k�3mZ��I�Ii��$O|�Uˋ�k���Π�XS��G�!��}A���u�}-P���{�/[4Mu�<�,�-�21c�?p��hS0�f�� @�G{�$qO��>Jgyُ=ia�����.@a9��P��QZ{Π��\	"/� Dn�V�=(���@_���,1�,����k|s`�-�#��>�"b��SaoFOc��b}��/���Ye��;��lZ$6�,�"�6A��FLߴk,��6D'����-5�_o�.���1��X��Ae��r�����]Rf�2�@4L��(�{N�N��d���2=�K-k5xr�����@L�;\Q'��BR&�F#\��B�-�u�:6x1c�Pk|�5J��pk������N�`��c���0�j�y�=���I�#Y���U��K'�.��2S%W��h��g�_�/su�4ފnf+L��T�
�hC���G_�n��`�8Q����8��%W�'Y�PID��D7!?պ�+S�����	u����Sq�;z�/���#�����0?ps�햫L�ٜ�3�1��̭�H��������ZNV������Kq���EU%SH��Ѣ2�R��v.y!���K�{@W�� �g�����S��5�,�b4�X2�-`,�R��'d��D����۹�ݺ������j����m�9C͵�f�K�*�tO��η�9E(`Kм�nG��Ӹ�w�	@UK5���E���E=�%�5?��#���#V��j%Q����<��uջ���T�-Ǯ�?b�v`�Fߝo����9����[xd��ײ
�Y��&]��6+��4��G}\���J4�=IQ��[��M�䡅��_$ڨ������k&�0]���u�͟X�u%�0�!�����i\W0��'�!Kv���[�x�JD�s//2�u2 N{�Lk�n�A��޲�1/�4��F�ߖZ��'\�I��H!�!�t�@�꧈��s8﷓�g�n�F�'���A~�E� �g� �`L���gc!u��M�,>���g�<���M���U�_���mm�äW�
�K��҆���AȜ�v��a�imQ �"����\о���A�?����n	}�n�r��/�P�����=��*�@��W$�
D�m;�(�L#ځ�GLM�W=ԋ�HOe����⥩W7D����nˤ���K���L?����~׺��~��I�+i�L���/^�?�� v��5taV5����� �qKQ^�sT͋��9���<g�{X���)ߛ&!��)��<�<s����~h\��bAn��Zچq�Gj�r��|�6�t�ʥ~�G��������E}��r&A֡��_�#��> ���W�L��nI��٤ws����&�kD�����3账�F�F��D�Հfdѧ@Z���Ԣr���_ z��ʅe�E���]�@�����鋏-�i%�VD�����L�|���ЧϨ#t��_��d^��SX�/�U����T�:5۪�s�v�J[ηUx�q���ѧ>����x�ӫS>�3���o�p�����M������$<1���*>ʬ�n�ō�ü�'��3\�F�RS<O�LCA�Fw�.����U^A���2K�~�{�|�����j�L}�d#r��K��*�պ��qU�c�(�k�+:}�{�g�p���"�����z�	��?�8 n$^#;�|do%����2�`�5N3N�h�
B�7D.E�����SnY<�l�Ej�4���Fl�.���1�ݫn�:���]��,b<����E���LA=���f~
���%����g��4��zmDͪ��?S�<�L�-�qKɔ��)�6�����iS��粝!ڞ����y��j�Ƨ�g����;��Sk#�&��bKc3�x�����֕>�r��r6�OMUoix���#����l���ɝV���|&�Cﱕ�-�;E��P�mt���Z��[�-(��L���4[u�+�y�8f GE�_r��ւ�.�T����Gc��N]��Of| & X_1��`�xsK_�8�+���� �u��CL^]{���g\j^�ĩ���dH���\~��N-���!�r1�t�_�?���B�R�]d�ܙ��Ng�Cm�XmP-`�N���|P��&t)�On|�/��cҔ���Ӎ �t7�V��p����GS�3*5���n�s�K\���Q���m��v��_�T�W0��1�Ố�[�}4�᩟|���iCG���7-�eN>����!��C�Nb/:�'�bP���U$��p9�0��c�%Ŋ,��[��e�]ׇ�< �ၖ �����D��?�5�f��q�b h.��4A�s�H��=}�o].������D��[���sV��.��el��G4Y���QC��%zjሯ�b-M|�2���@c��QQ*�qWjY��Kvm
��2W\Tr��p�'�|3ϗU����n+�K�x���gr����'�k��M$�,-��"_SpsmlD�~=_�1��b��_3�R@ �CǇ�I'����l�@G�Gr�w��a�o�P�f��S���S&	��x�����˲iCI���/r�v����t�~���-��=����p��+/�U���/���\�X��0�M�^��`g_v��C��e6���8tadV+Ø�-#�qY��Pv󊮨emn���!%�Ͷ��n�������0��mk���-�t}?$6����G�V*�~���T����{}3��3��s96Ĕ�ÆD;9�'����Z���5�C�����CQ����ݷ��!� ̬����iphXX>%˧��)�;Ns�o�}Y!����I�dn6n��M�;����Ɲ�{�%E�?RK��B^�Ȋ�{�S��'	&�C�[���j9e�!Opp�����Pb����_"C��)�z�g(�Ė0URn�`��4��=��o��bX!~i�lOc����zO6hE��/���b⮆�CJ�}��nW:���0�q�� ��F�
��X��*R���+��;�]m���	�L����/���yŲ�x0��;||�?s��{e�FO�����B�v&�JA��ji��L����|׃Ľק1�SD�� ��vO�H���i(�Z.X��?�!
J�����"[�3YXБ�)���`�r?wP�,�p2�bBxMCʡⴐ��K�TZ!���[�ǉ���g�?�/����7l&u��]ײ�R��[�=h����ؤ�Mj,�<����e*�L���v�@�ٍ#P�f3�b���q���6��* ��IB�r�]B���9ѭC������tZ��n{\���53!�`���l%�-��	;(/<�q��R���?�1 �H�����d>����o*��u��r\�p�T�X6��G��Q�h��:�}{����S����I7��T�m�C=f5��ޟ�1!q!5>o�w�Y{���w+6�3�%�T~�o��ʑ�w�ς��Qg���6B-5a��?D����P�Q��nh�Kk%�Q�$���2}1P����>9��9�o�:�ک�a�F>�^�z��%�9eVf��k�8$��S�s�"���rEي����D20"�ׁd��_���%�o2{�}A/ۤm5ԫ��ْ�̭c]�G�;�	�GX �� �V?`WC�<d_r�*��Y�N�m�W-<�#�>�Iw��+^����a�+0?_�u�3I �v"��B�B��[`��4Gb���t���V�d�w��K��/����R6˟�P�\�b�b�>,�l=.]�$*n\Q��U�u����l˃Z�ܸ�[~����t,Y���*�������0�k(D���Ƴ^ϲd�■�uXYt��aH�=�}şޏ���do������I�WY�^K"�s4⋴��!� E�[Iz-���$&��B٨�[�GD���Z��U��p�Pn� #|닭T+�_ꕼ�����Zj�t8���R���$n��[ټ���6t
��/ah�����<[O��0aZ�'�H�+D�t[�@X^��Ǽ#e^���r=�%Q��A!�<+f`o!f��Å){�$�
�c��A��ݠ�ȝ�!G~�/qdu
k������|�T��m�[C�HSH*=��:�(XL���%DE�_��S`��,�]{��à���BK:`�$����ҥ�0g�\GA���ۥ�T��?�CȜ��2��X�L���b_Z%�+}����a����WSf1�h�w���<M"J��g��p����Y�xϸ��λD�V���5��!��b�>����B�}Z���wa���K�JN��]�%�:�U�8�x��A���)y��>"(VU�c�R�|%r���C�����V�ԣe>���c���6�6MQ�{7i��+o�P�������j�z�.\�Y)� �N�6�vI�d��_�p�6ɕ���Кa@�[��9w�����w�y&�ۑr�m*�>��*20��U�t��z�o�:	��m�����^����9��{'u�|'�+"m�{ ˌ=�y��]��
V�c�2NKiR2h���̶*�V�����F(����0v������F�U;��Ϻ����ƵQ[Z���$6�"��v�'���$�kη�W��F\��gU���̲�=�,�EG���ĉ~��r�Bp�N,kQ��A*;9<D���i�K=�9�*Q��ňc��^���m�x6��σD��a!�\�pT/r���&��s����[Lp��'=�/}P;�����V�VWXP,g����� W�F�%j�Bz���-pr'��ꁿ���k>&�D�30���-�,��i��A��V�[ oo� �t7wR7���_4��Fls�9�q"ς��mxDU�GUd2[�4�ӎ[+�T�\�p�Ł �f�F�C�Ί3�h��_�֛���ge�!�3e�������ɱ��ѐ������k�[k#��yd�cv� /����4%!w�~�F@E���M���j��S��m�N��>�E�qNn�6yi�\�����c�B�~�}%	8ה������'���qϾ}�N˽EϜm��']B�����070�S�IA;�fe���e�7t�7���U��#gT�矌"`N��qd����v���qw���H����%T3-G�>o�sˈ���.�/��)_�
[nMɉ�;STcN�5ku�����@�P4�
$����rn^�w6��T�	�aCu���4���U* ��:�ؔ���G)�W�V��>�����5 &�	
��8t7�$�׶T96��UC5v��ui�`HŢ�`��5�:�x��3̧J�^r������)���nբ�r�W贈�Ms1�swu����k�� �Zh�%�����$"�އ��<[E�k�4[�	��r��ㆻ�~H���
wJ͋5.�nlyY� ��9Ү��o?i��n��m�����n�I����
5��3.7)�&Y���Mb�Pک��/��lc��%2z��^��=2.G��@����&�v=�ǹN����֥���K-?��y.ߎn�p,�� v�����r�L��:K����&n�^�nu�]/ϝ�s�.�T�Eav=�4tm\2:���k��}��oQ�mn��d;�p5l��Z |�1"�]3l	������-l5zF�i"�Y%���CO�l	a;>*�>���`O�JE�7��1���ѧ?�{=-�2v[����Ȥʍjz���u $�{��{��
�'o��D]�<N�'c�������w�
���yFU�3�U0��<��T'VS�X�2w^�T[b�ܬ��]�'ܔ�q��!��Vd]�C@ɯFt5
Ц[+Q�ذ$l��畛�rd�$c�'�ҕd�%D���4�|'��y~$��:�c�ȷ���S�	ݮDr��GDN\�.��I�;JЧ@<>ȣ�N��_�D�FpU����-�����g��v�5\u[�0wYU�;"4����$�N~��-�H���ɭ\�4��mBeh���1V���P+C^��O�ʮ i���b�	M#<�e���(_%�֝�iJo�t�����x	2�L�x����]�эia�\k��in�,�+F�ba�w Zn��}5*b7`-d��l���wB9�Bj�C�>�p=f
]*�9����f:�TS6��u|�ɚ
x��� ��J]f����:���Y�?�[O\xYl�^�
�pCAwG�<ğ\��/Td�g���3��7o�pb��A�9xR@���<�����E��؆ �D��Q�Z�"�댕o�xF��Du:p�ĺ�3)M���+�z9�hF6<�)$7�cF�����J�+Y�/&t��4���2������>R6�ʢ�0����+�������8�]5<�k#��}A��w���N��z@KO�埇d'���Y��Ƒm�?M�b�f6Ҷ�U�?	]��(c��h���k?�����=�%��wu��:%�GQ~�ա��^���ȑIh��p4���'��+.�r��8�6�6z�O�T��L�)nmpB���3f!`k.�-G�/K���N�}T@�[���9ݷ�������L�1��īl���t��}��f��i��A>�����g��0�Mp��d�E٦��\J����������4Ai�	���KmI�}8���dG^(^����F| ���.zUU;r;�A��g
��xi��H՗�||���Nx$DxN��"�އZTާ������@�c@?؁N�����W��!�/���Yhr΍���QcQ D<'�]�9��pil�i��]oa����N)���"8�ZM�ѡ�@ E�{�2�4���/��@�#�"�˦��-�NX�6�ۗ���nq����g-��R��Dz��^���Q4�Ø�(��1���_�j���^��+.ʵ��x�F�%d?���N��6�`���Ԙ�*�o�Q�k"(�1 !t����2H��t�<b2ŊBf_���pN7�b�$Qk���V
Y��wmI�ۣ�:@j����r:�}W���Cc�[�8\�a�A���M�nXgFK��-�#�Bq�%����]y]g�Pj{7��T7��kR��t'�ad�|���8`�^�e��7�(�|<�i�P�|��3���R��%z����O68�5���N"H����C��t� ����χ�A��5ǧ=Mf�+o���#
�D��^������E��^mT�e|=<��fl�asI�qɧ�s�}��)����9ʕ���~)�On��vj�
֍d����g��$������(��!:��#Rh�Ph� �7B��|��!�(Iw ^g�a��̢ ,8E�L,0m.2�v���p��A��4�#,�ǞG{��>� ߌd��-݅�=
E��u%��oKC���D��Vp�Ik�>�?�r&\�Y�2�}w-][�M�c� � RvE�D��d�����OqF?�>:<_�z�I�HX;�Qge�;>����%7N�O�#��M�1y;I�d6���#`�Q�Q��Mn�+b�"D'"��>�u�^:bRLX㣠gz���B?�s��d��|9�E��cq��a2̹�rH5}*�q��@;��6?'�1�]�)���:�P/�j��ّ��Jφ�s�G�[BB�5߻�x2�1Z�Jq��. ����j�l��Pݞ�Ϸć�/I-F�Qzg���v��a�@���k��Wr���3�>L��[;��2�*���I 5cl=�����ڱ�,�H��W]��Q���.}���/���o;[5���o�7F��=DÕɱ�	��}�FT��������թ�m�b�'��0MVЌ\y�����dr+��'�2T�%���'I�.m��OPad�X�g'N�&�/����.<t@n
�o��K��B�/T3j�L��e�fo.���K��ɞ�k:QyJ�Q��"F&��vۇ�aM���!�+������z�>cl�`����}r���g��'�����������S>�^��mOw��{
T��!f�&n� �w��;,(�r,�{@V-7CZ�ܖYQ��[2|:s�e��
�f�4��L_��>��5�P��/���n�Ĝ,�{- R9���ma�*�:bWcQ�	&5i�!�,4'��]�����#���SQ�K��U� ���S�lZi���꭮����c3�_?�P�V�� �\����O	B���!N^����k���ZŊLBّ�ԤK�[�#�ebP�s���ybŝ��9!&��5����$l�F�g�{&����=z�#�����GPE���(���^��c5)S6�8�s���F��3�bL��m,�1����v1^��vk[y(tؤK}L Xw�t��[!~�%���R��$�����;"]����Q������Ǔ�}~l	Tڗ�L�(�\��n�)gb呾�vDQ��c�[/�g�0��e���U��씉�(��5Ή�'���c78Tvڽ�B~�4��XgWr��dݭS�!R�_ ��b�_^J����F���`��� ��;*=��Ѵ
��|����j:��tJP�����T��
X�1H+u]CV߀� �2�*�9�������h�b�C�y2hq�o�>Uũ-}�έ�+��4A��$Q�!�<�%cc]��2B+΄� S����p�fN"B5-Q�v(ErN�e.����}�*�e!,Y�=�$$�Lۧ�w���/j硙,_?��?��@z�6<T�(b'��=�~A:����1�8���qaY�ntTw�|rP���d���խ��9_�����82e�*���o1=�_+E�-�Z�Q��K@�*�4�&C��, �%Y�����1?j�Gp�T��8(@����8up�|Os�
��W'��H�����"F�B�K�y@�o�.bb�^����qBe�1�лq�p� �}�>�^�K��m��a����򓋏 X��t��V���R}�r&�E�X�?'�50H�R�H�O"}�*>ë�g{9�H�r]�oc�`�[�щU;��Im_�� _��7��W��K����h �Q��U��΂dx9�	���8���|� qD��.e
�汩��f��*�����!� V&�(�J><`�L劲��xo�h���$���5B�a�@�c�t���
��6I�&��z��0L�ɝ8x��ư@�d|9r��:�%Ui��Iݦk�[mƯ�{E�C/��c3U��S�?
��r�kCj��xMkR��t�^H��I���� 7?��mxSG�ax��d#�:K�d[�Һ[��ґXԥ����8$��קgQ�a�0-��U��Q�W�9怉Q[��ց��S)�Ҋ���\H�Ĭ��j̈́֜���S.�ɔ��,�
T�"���u9��Ⱦ�
�ၙJ�l7��Ԉ��'���O���3%�י<��f���������+o5�eo	*�?��o��`Q�a�>G_Ze;@���(3�ʥ7��e�:���[�2T���'�w�T�Ff�����$���."�.�j�t�˽��)\.�a>��rޔ���P���cB�6��pyB��\�g0��A�B#�|��m����=t��xg�X/ŀӏ�y
F��6�TW�@�*s�xb�c8oq�l�_,N�0**Ի5|ϗ�h@cf,�m�JAe-S�5���i@��ZL��J��Pl�P�����B�L+)D8ū`<�	} n*Pz�nsvQ?
e��gs(�ލ�	�οoAo�%"*�FN;ka?ܕȋ1_@��HE�Xzd����7Ø}�{�&��~Q�|1�&��/� 1}a����2�\=Ω�(Gt�;?$�'���4V;����r".�(����d#��/v�|1Ui_�@�2�V�V��� �� ���%Q�3��T�t���Г�{�����$����\�Lf�h��YBQ�V�kP�E�Aߪ"J[[��ԂzYev�H���{���4��-��6Ypk�Q�Ev�u�y�z�g3&�/	ˎ���ܹ�r���-T��Q�u?�Su(A�o��*P�Q��������a��ƹ����_R��a��gt��h���ݝ���D�2"�� t��=��bx�a}��jp�ֹ��ğ)_r`��262p�ع�Q��	R����@i����l���.\k���A~eKCt�M%ۏo����2��r�x*�<��k�#Eܣ���nM��P�%c��7���S�@�'���w/{��T���!� ���f��d��mjǶ��~lʦ����fU�g���E�纄�]����֮�cq�� �qS�B��s�)��H�)1ɔ	�Z�=�Z�z����B�{��8����-8�g�;|��9�Dy�e���q��x�1�Δi���-ċ�l�*�r)ߵ�s�~��۔�^Zf95���3��JAX���Uz�5]86�lC��I 8I��j�q���m�{���J�9"Q�B���Q��Sg�����y|�q�gS#�SpV�M��~j���Q�RQ�(R7�b�|h]vU@L�wƸ��e=���M�k*2�/]Bv�z	ר��&@~lHE��װ���٤a��k@֩���2��+Si�Q
F�M�&[�'�A��M6�����$Qs<��PH����%���Aq3����I���]]ݚ�A���[
�Ͱ��p���ΙyH��s���\s��=��c���p�! ��� ��H��7����R�Z�����rx(�f��?L.
�e�@��Y��䨘�IM�u\�P��S}VƩ���b��DD��M�󧎼U��>gDmd@���r��o�D�64 :��dr�.�� ?���ń<v�w���N+���pI�L�OK��d�k�E��P�o�'��+����-�5/�M�e�4����Jz�`���Gʺ8�L�]�@R*��2
"1/س�D�{��@��4-�V�lȒ\D���7*[�%��n�E5EWf��"�f?�,.�f�,˝�X�7��_?�W����Qy�ϏG�C�Pf�Hv�(���%�#�.U�w$D�e��_�>#��纴�P嘥V�i��(�o�p���1'���E���Wa�K��u:Q3��Ξ�๵�{�I$��!XߝT!�(�i�~�H%iCi����3��
΄��ٟ�K�\�/����z���*�/n0�B_���ɑ����8�|�W8����0�,�\�x�?��J���&ǔ%�q� m��N��}�O�k�qS��L�p��𿖷����*���u�H��G��B'n:P��؀�
��ɺ6мL���R����|l{�(
�6}����4rס+S��I�3�����d������z����_��e�)�(�s�����o�,7�2K���<P�N``�<����h��+E�'zL	�?��5D�|��tc:�.�_սn�ݍCF��ħ>q �97R��z�nh��@�Z�"y5M��4�\�߱-Dא|={4�]G�����s�"�8S�H�lx.	F)j{w�=7�m���2*�B�qą����y6-��F#���-]O�M��$ֈs��?,t�Gm���Л���:,��8-�㓍�N�T�R��0�EHr�w�5�M����JC1����̽�b�ɰs��t���;"g��E�Y9�}HtcU:���Bd�k/*~�Vj�L�#Ġ����k_�G~ꆈ|FT�������+���֒�\-#�^z�%2��j���n�μ%B�|x���;$^ʁuxǇB�Q#�|���ãb�~"��E h��gۘ߮���n�:�[�e.jgf���Kw�o����5��+(�˨��6z�����s���6�"r�H�K������4?�jI	��D�>��񂞱�'�~��=r�dbwQ
�2�b���AFEK�̱YKj�<���~N�^a�$+
��]���{���hGp˓M��ю7��{jf͑�ˍ]����_��B�l�t#e�PGU�r\������C�9����t�:+
�/"�M��@���3^���v�e�O(�Ť��y��ebfQ�>֟�ς@�,���u�C�D@-��˯HF09?G�NO=����"'��ٝ�7�M?פ)���ˊ��?���:T�f����p,;�ogua��p�����[yN�1i��˱%��fh�,�*�^ܺ�6c��T�WGЊV�}�*<�se?�f���O�	���x3%��zZ���6�^�l��=&���S7����G�qS���1c�&E������H�l"����w�M*�q����	L��z$
�=D�ԥ���b�+�q��ʇ������5]��-�g�r�`��u���P����������Ƽ��*i
�t9�fޢ�0�,����u�����
)��{�k�	)��\�R���ަO�������Ƭ�Xc��$G���]���w{�Q_�@����1������) �AV$}��?�i�^���X����:q�EK�`m�;�ռ3��o�y���4��i��c��b*�Y6bU��a���mI�-dv��<+�|�y�f-@�3d#�a��׬�J��/�7B�~2��v��Hvt�)���̈Ur�a�å��i[��VK����l��w��M�7�Z;e�5��[��"]m���rA������d<�5+���ۗ�̝n������o}t�r��b���}�x�;}�a)�M=# �P X�&)��'�qirM�`��Jf;#bҳ1�������S-�`eUt���&g�>~~�y<����R���b��2Xϼy�[e����j>2�H'��N�Q#Q0��@�;�K�`�Ӟ$�t��g����/�Q1�zUM�+t9qB�z�}6�����u�ie�~�"P9��.�5M�@,;\] ��S釅�R%�'��-�����
z�`9�Fj-РA���jF�Y�j;�A�i5f۱�R��~�ܹ��:�4�5#l34x���rOF�X(~�E���΋�Pke}iA�
_��ÓH�箦]D(�\;����*�2JT:z7�L�"y�r� ψp�3��H$�����y�Cdx�g�s	}�TGD���_������%,���,�畆к�lF��ui�>nQ
43n�n��L��ލ"����cb��BF�y�1�z	8җ����������pW�^T^!,Q��ǚԵ�S���0v��w�~�3k���ɧOD_4�@4�=�B������H�X����b�<Ջ�Voa��f���n�X%eʕ���rW�0�ۻ�����.
��	�C
Z�ʃ��ΚB�P�m�K�Ym">�/��Ec��ޣ{Kyjx���t�
�Y�-Z����'ά�:�ǉ����!��+��z�c�t�v|��P���IW�m<v_5A�����d߅ڮ.��:�}�x-Vh�b���d��yú=����E���'�u_]�c�v B�5yÔ�}!��ߘ��U��B�3)iP}
�G��cz��"a,�n�V;縙�N!W0h5g �or�4�9橪]O�B������a�+�o���	+�H��z�E���zS� 4˗{��
��!�n�X��Sr>-hPoo.s{ș/�_+�}��E���X��砋~6�ɷ��⯔��'Ų̤��;��e9�L����������ʢ�>��?�@��K���B�[sq�sz䉁];l�	��C6��4_v|��`C'�r��Z���;�~��*�XA�e��m䌧�c��Ds�WA�A��/f�J�X�kQ����_L���MzR�Vf�>.�4ׯ�� Ex+-��Q�	Y�ʩum�v�vB�é��sW�DjN�o�e�w*s��b�K�ǔ�xU
M�]�����v/��8_�.�����(�kI䙩w����O1�X̶�4��M�0j�w �Eh�lB���J�g�弙u<Z�5� ���UPCG>a1�_O	D&�ԟF��¥����������Ƃ���_�����N��Hnr>�[d�a���)z��d�lN�dqK4�>S�V����`u�"���*^�pw%e����Ѽ�P�RC��?M���'G�<��4��L �0(����s�ll�8'�Lu�`ta��"��@v#aLtu��U%9qA�
�m�/���Ք1֏�������ۅ���m�����}��]�
z��U�K������.����6��FD,bBQ6�4e���Jΐ�s������q���2ل��6:��ȳ��5�¢���t�h̪�4���})�~]��5��O�@���q'�V�W��d .�c�1��[��,�$%��uW�-�-3��/pjŇG��_S�P��2h��l_������2�{����;�AŇ�7	����3֫:0���&O�{�Fʜ,�Zu�_��0�10�-���OU�7���`���ʤ{P94�W����O�@��������@q]��v�؈��%�/�c��W��~��+a8)8+������>-X���#�y�b,?�k�#�<eҦbrxp̢���ZT����=rKϴ�g��%!�5W ��o7��1���b����  q�C�K��E� �IXF��xw����J�A�\�~�e�j9x2Z��>���rj������,.��N�zn���!�nuU�)����zC�놻݉)��@Zn�?JLRwk�Qd�HI��T7��k�0�D��*,8����AV�c2�t|����H���YP}�}�~�5Am�~VK��=��o ~��2���X�� \m��22Tpa1��Y��}8mw���|_r`S\`u'@�/t���IR�{����T��}��n�wkVB�L��קr�c��4+n���Td�?c��&���$sJ����KͶ��$�祺Dd� ĵ��ԯD�JEJ@����j���ڹ��մ�wq��9�3ζZ�J����ܞuJ�q��r$��'�S��a?:A�{x팫�e���� �E��
�T�e5w�LV�KFW��Y��J>����H_���m�f7>1��V���H�t����JV��Ta�_i��9�d���7��2�a���7)	�!V6c��P��*B�xv�#�8��s]��'ꀪQ5��Þ�}�'��}�������������XR�|�������������a����P!Η��Uz"�;&j�V�#�|�������������{� ���3�h�x��u-���lO�;�%`դp�3�Tv=��*)��)���E+�^��{Lm��.R'��x=oy�i�"��0yB�l���b��ӎ/l�?��)v���}l"Yԡ>Q�Lq"jlťi�\�ez�,�0�$%��Јw�>�[h��a�E�-' �tM�����#=Lif�x8`��z�I:�>H�+>��꿗��!t��Z����^�c�|5`�*��bW�pٌ�
���v���P��pl?�|��IP}��o���~N���+�q��g��o��m\nA�`f�ƣ�}���Z'}�0��\�'�ʰ��|���K����c�#����V�����ih�9�f��NM�|�A���z�p��.�S-�p��03}A�S�
-}8�%���8��R�yX�8 y������9F{O![o�q��+N��bjܣ��
�E�&��uث�\���;±���U#@|&�𶆥d㼊�#�C��[BqM�di(Y�����ꤘ��mm�;����e��PB��c�{��T��J*�y��S�E^��qj���A�����ko�7*jr	+B��i�.��:�<�}i�w�!���!�=R�t}F�Wao��i�8N��~#�����N�J�3j��=�[�ȸ,� �c��m�ۋ�`�b���TE��kzi!/2SF�1��n�	�GI=�i�Cnu��,�ΏBf?��p�F��SN��0ں�7�L6��~55���\�
E#a�v��?i̽JˬV�񯨭���X�e"�����K��[�[0���fҦ��H���L�a�{��ќJ��ʥI��������lܟ�2jw,GL79�(��:L[<��彉���ޖ�)�xwvJ��y�� Յ����ԁ���1\O��nT!ظ�~sV0$|�Ÿ��ޮ7�۰�v\5A�Q��f��u�9����<C#6V�۾�J�<DLm���,ɚ� ��v=mp;�PgC5����7�E6t�>멈�'l���q�ˤ�����&qE2�����I+b��x�%1~��� �����&��p{`dc�w��҃���A2k�Y���E�e�f�x�R~}(D��0dyl�E��w���n�sy<B9!e*��n��_^��K��BoP�f\��b�3�p���T�
"U�ptZU*�����#D�H& *|^�&0����_��q�ʤ$T�}�������g� ����|�S��/*�UO���v�%m���
R�|d�����t�26�����F��A��(*#��u��mʟ�8A�����ׄҬ8Т��ߔ���-@�W}��1�����1�B"���<2O��V�K@ǣ����������1H�.��H;-l�݊�m�?�7���z���*&����BZ�}�۸��A�W#%�rC\ɬ�8~�'�`�߿�;J�s	�1��O4��a+wB�}*lB[��� ��"$e�\:y9����q�j��8�vUd
A*j59��l��Jq݋�K�Qd�&�:�ȋ�����[������J����
�O�4R�Ҳ��ЂB5�-j��6��"5��*h�F�4�9g_���&;.�u�_3: �5�ѥ���ϭݓ���� W����;��!����˔��_�� ��{��G!�e�j���!�#�:=(�ʑ�zV�]h"J�*>�͹P<�-q��^1��qp8������U���~��c���LXO�^W0���섖��;]~Og��L��Pk#q.����r�5�q\øٷ=.P���_px��I�5	�^1��T)�҆|��g�LH8$����7���Wv��C�`��T���l0q���B��'�����~���G+�+JW1��������.5�X~Ļ�x�v�T"(yX,����F�^ ��j��1��Qc0@�GIw�\K�`��d�v-���Y��`��a������(����Y��G�ۤ<���4��,2�����U�:�v���8�e0ys��L䲚f��E�n��+x������й�����bʂ:̣�/.=�lJf7`���ƫ�f�B����Q��z�f:\��LB61*��@fɜ:��x�7[�Rd#����3��
/ھW-:�;mI�����E�v��		Z�IXp�Ǭ,��+�;����#�|��.�5����F��ki�&�������d�i��z�������)HR^\�-�d�{�@s"͞�Q%��`�3��Ks�P5�>��5Ut�ޛ�@�#�M�u�X�埆M�8Nk
��" ~?)�V����2L�I���a�Rq��:C��ѹ~�[��Ų�m�Xg�V�,�Y�
e<ᚒ7?���}5,�C{d"Y��70�BE![�d~�l\�"����ѵs2��(��8���[v��ԟ42B�$��^�[{.FJ�1�����E�Ah
3��%Eh�����n	+�)�i˥�FTAO�V%�j�9l��""i�H�jK)�Ө�߉ Dx�u�m�LY�ݱ2h�,�p"K��� ��{!��ը��S�t�X�^���1s�(���`����EQ\;��5�����=��&T�]����+�t�9�Lċ��������n��BqpNnʈ�<=�yF��7-"��p��������fl�#��LM��Oϛ����yI�W�����\ ��C�w�x�P!�8qS�p�x���Ĺq�4�&�>��o�g6��Iz�'��O�a�62�971��V��+<�w�Q*�C�lVW���4��bar�|:���ġ,������E�J)� �Q�[�p�y"��a��{�z>��kD!y�U�!
w��Q�(	�$�5G�<'Z�G8��q�Pn{hFx>��tJ�� /�	/P�@#�{@y���P������H��(��J�����+a��Gr +��@:H�n�%A�x�r���VJ���[ޟk>�H�^��I+���Ԍ���o.�I����Q:vk� ��ã�{�7�q�A�F�q�i�sI�p���e�C���j03����'��C���=�Y�,�%��>��n*4�[\�f�/EY��8}=������.��[�E�t��Z/���G�w~��Ɩ���6_�������� ��<�qM�`X��\QK���y���#�n0�˃��}���)�;'�����k�N�.T �VQ���<p
�DH�ID)���}�%/u�&t�*���Ey�;eP��gD��J�B����r0*�$����iY����Aķ�mLS�hѵ3�:�a�����]P�T��,^�Kֽ�UU�������榘�T܂K�~�-��Ȫ}KޛrY�6�:�ikM����'�67�'�"�^�$qe�������Q�.�����"~/={��S]xp	�u����&�wN��b�����{~n�_��@�	�wA�(j��І[�n�|�%�W����]
�s����]�cq�%,����	��8Sz����>+'q�\�h�(��Q�~���~p���2��ɥ+Q��5�a#���yzA�Z�qcO�t$3M�£j�YP���G� �ᤎĆ�3���ʫB'���-d,�sIbT�/��9�
�9=a%��%2��Q����v�_OU��gW�v�0߳i����(�8ՀP���J���m�b���+�J�:1�K���rN+o^4��W��ڍࡥ1�`�[���C(m1lK�E��b�Q������3ʅd�d͆2���<v[R��O";����v��]�o�a���v'�h��P<	&���ܮ^Y�e�l&���Cywf�xQ���e�
��\�.�G��)�+��#�'8�ܻk���_�R�h�����9�n�Jw�6=�},H�ة-�p`�?�wl[�H����#���h��@�e�;�*�D��נ��f7�#&X<^/nˈ���N�+�8:��1�o�եds�)�8�&{�����sG�($�׎�'�u۔�ך�l��p�P�5��&��ozsCLs�9R��6婟zcII{QU4,��<p�^�kg���Y�����m���$�0=�	'�5w2#���07/py��;�D �9�J�U�� <�QD�IVdBǛ 6����T�IO7Z!����Y������~?%s��c�D7��T��"�|�$W�Yѷ����W�&�c�͊���+�ӟ�?K�Kq`��ȳd~�/�}_�链�k˔�^ٜ��Q���e�"�Oڟ-1�7D�I����Hsg/�A��(� �F�Z�g��D�9I'�\�[�ؾ�(���]J�����hc� ��W��dt�q�XGDz��=��ĝpQm��
�=�YUSD>�<J%~�If�cr�M�4��q6�{3�=��k4��N6)@�'�c_���L��aKL����IV9	%IԠT������Ԧw���H4�}��j�)[c�����d�x�ɻ��X��P�"5����{"#�}��a]'�ג˄?_��J�Ȕ��\�rS���K^�ϣ��v�ǌ<7�"k�u`T�S�F|+�\G��Pw��(���ֺ�e�eϙ�\@ �We����gr@���N�r�:|�6�Ş�{n�F������
a2|'�AeQq�U��Q-��Rj8�̭dOJ|���H��Q�������:�`j�W��W��$t�4����w Ф>��u&���<�]l'd�V�]��F*�@;)ejeV�3�?��k����� ��V,�^o�k�0$:�S5!�Fy��s�s!��t��N��q��.�\�f��D�`��rU�BQ�|S�K!h`
"��Wy��%�Ա��r���Gz �t�����h����D��� ۰&3��)�>1->�-���-��<�Y�5S�S�^��?%���M�����9u<�2����H��tcHB|H��be��� d)3H�P�KFn��p"��u�P
�e�����Y����74�+��	������C|�eAǧ��#��&��önwŧB NPy3~����������������F=�wG���w��@���Ҥ,	޳�k3F�K�J�9%��˝��2�-��������Ob�$=�7����G�+�v��!���ҹ�c��$v��V�8|3`�<&�4��4�*��hQ��@'A%,W�����&
��6�ڽg��ca��5��Edu�8!r�x쟝�N�=�R���]�%`8ЃX���yf�~�i�T8�%<�5�C���Y:,
�ъ�f��,:)��Lb�E�f�����Ml��h��B>�����M#�-�dzqJ���Sζ�_�
 oj�1)y�4�g
��,Cuu)Cc�!ϼu�5�ʦ�rժ����d�w�`�u%	���r��D�dx��v$;�����Q]����o��P��-�yK�l�5���3KV^����qX���g����p^^�AQ-T )D���Q�j��>$�7�#�(�TVX�h��NnN��"9�
�� �.��y� u3ؕ,q]V����p":Gꖗ�(�1$��z�M6ט<�eC0��7玞�/(��]�t����$����|U9��*x4"R��1�0���<.�����c���J+�Hg>E�!�����D���[���JNA_�7[�L8j*��s� �N�����>꼜VN�fH|C\��$���WM�!�/A��
6���܌u�k�R��=A!�hl�Cg�W�u��?��%ׯ�8f��{cL|�i��_;J5���p��n=��U�7D����r�=.��mN�F���1�?W{ֳ��¤�ة~��㓙��V���:�;G�F�0�wG�y��KL)EC7���h��Z�D<l�:@���T�����$�9o��NE��!%('Y���6�H�i֣�W��0�9�`���ϥ�M]�PD���Y͘Sy�'k��V��Գ�m��&�H�<R-c���Ǚ{�~�Y�)t���ۓǭUۖ.�
��Ĝ�r��5��L9ۅ�԰��@m�l�����J�rn��ʻn�/�����k�~ 1� ����~�M�6-FO;��z�rB?���Sk�;�S'�j��	$�AD m�q� �/�q�	��G}�����θ呠�g�e	�= �b�N��u#I/\+��	�;�c��U0~��!�:}{�yq�I�� ƗG�vo�C�Mj�!`I���0S�(*�4>��m�xa�>�45Yt_�W�ND��rӻ���u�xJR'y��Bp�w���9�a�>���Si�4�]�m"�)�w	��k�m�pj9�2r��������~v��/�jX��'OB/ �Ĝr4���՜���Ӈ�~%��1��}�|ٞ��C����BT���֯��ho
g�3Rf���+������l�Dխ 505T��q�-����Nh�v��\f�}��E���ߜЀQW����(j ��.@����z�|�7ǖ�������~�/p)X�ǞH�� ���k��3|�I��������R��h���	v/*6Ck�u.q9��"��Z�:-u21V���1�C�q/��I�s�T�|�������h)D�x��켾���E:ǉ��N���v��W��Ԧ�䞦BK� @]�/�]��ȷ��!Yx�R�9Z"���Y����k����K�fŶ�D'��G2���Sz|XH�ۄC^b�����Z�V��_��ؠ��=Q^�$�ɞl����@�.���#�"x���*�c�i�̡)�H�8a��b���m���J�V`}�����Ak;��"Ti����ݓ��L�Vxc�m`����S�� �V$��6#�F�9r�gx��G1�-��	�)�}���a=���zUΏ3�/�l��4�`�kd�Ĵ�%����2�`��$����4�4��~]�q�\u����Z�b�ډ��ߟ��Ҧ'�� y�m���3ǎ?�k�n�P`G�<m}!PAD�x5�|��\�\[<�c�-��	�+�7&|Qօ�0%mH�?zC�	}�s�'8�`®���i�a�C�8�$��M{&����6��=�ӭ	p�u�R������X��Ixp�>�о\؋���NLukZ���E�O�W����bY~�s�č�]O�g��vB�_��S����g܀�9q{�U�H}ܤלT�L��;�g����҅�cy��ԗ0�& ΂֨72��1W~֭���X����H�g�[�q	��j���u̦�����	�T���D!��&u�b��a%bF���p3�ˢPH�+x#C�����Ȼ+9۟��m[�t)N���X5�ŖRr���-�!�5��=�[��*��&��ܰpT����[���({�6	�8b�}N�S��]i���\�B���ک��R�0�q$+U%DJ�/F�Q���8$&< ��?^ϔ8��h�M�aG{�`��ف�kr�J՗˜Wu��~3�y�ܚY���(����VA�yN����9���V�P���o-v)�QH�*��쒉�}��4����X����*�M�L���&�����/�<�R�8\��2���4|y��<L۞ ��#�%UґSn&M�r�b�^
@$_
3&tԊ��?W�z���'Y�X��/�+�{k�="������s��J������MD��P2�R�Gs�zn���W
w;2���vȋG�9�[	��=�\���[��@����56��n ��9
~q*����aܹ._�W��C~v A��y{0}���^����zexc�K��z��\s�A q7l����ܣ5'�V:*8�:���t�'d=}�]p�5J�ƋK�S	�ĕ��T�j��V2�
vl�&C��X�3x����} �3z��6Dr&K�!nA�O6�Hc)�?�TxJ��!�E���4�!>$�aDext=��p+�5Ԣs��]���P�� N��N
��y�m�����@����_	�&��ӷ��;g�	��E!�4�R�g�DO�P�M�m2��g�8~~m%[(|���:49@�@Q���*��-XUM���CS�u�f�F&��]�vb���C�<جh&u�
������&�&�c��!q2�N��\���T���\^�N�n�ğ�Q�G��(Xt�7���E�ZU԰��wt���f�~7*	�j�9������Z� �̔�+h�Z�J������tÂ�Mb�\�Ip�~b/J����"rS;}�/y0bpܾ�Y�~��� �����R����2m$�xI����"fs(�3DD��/�,VD3�h��0Jlߧ
ط-���\��,^;�K��޳&��A6~�x�n�r����ÔR�T6����q��]���o��4:+s�&j�4������Ȭ�� ��Fe�d� �@'T���B$a��N��]º�l�ҬEg�����|�1�	�������
D��"f=�\V6�I&>�{�)mJEy�QU1��U��M�m=Q����hhB%}�G���a��X�>0�xw�dE/��FK
�����d�`\��B����ۧ���A���/���n�Η����4ܱ,U�@���9cI�W���d�͖��\`r�:��ƣ)���b�ׂx"�9��4�ܣn��o=}�n�OH�g�vTl��8�)H��i�������4��#_�+���_����)KGOD�l�+ٱ����n;�W� f�,�G\��9�j�dOu�z!3��jB�HgV~�j��k�4Mh�m�&�c��� :&}��:�Ƒ2�3?m1�������co4G
xw�3�T��Μ�&^�o�O���"u��Q��Φ?s�s�H�ip�q�9%�6r�y�}��_x29��%5�y˓����6�H{�]AFޣ�]��e@�rE�Z�W*�6	h���e�RW��:�Z4jUR��9c�(�W��Y�AG2�?���
��1�� �ޔ���"P|��Qm�p�\4�{��1y!��ox��\�� �!��Y^625;3j)ٵ�r�f"��t_2�i-at��8Է9j�$d5�t�����BA������\��@:�3*}�O��m^��v42��rj�L�w��g��2f�Y�/w5�^����+
�|�wg�`�A��w��!:�M5�,�ԛ��8���휺��Y�id�����W"}l�W_󡓹���xG�\�^=n�]D.��貇���u��Tp�h��Nt�ݯ��3^�<އ��	Li�c/.�����C��?_�'/\1`�#�^�ٱf#̸K퍃��T�=�@�i랢�+3H�\�h��P��I7�� [�L�6υ詠з�i����?���C%�a�a�//g0��K<�&�HbO[e
����f��)��u��_���V�~H��bm�F�tR�=Ny�t���ے������ܭ���_�����l�F��[{!����[~��di/����b��oQ��,B�V농�o��mE;`2�-���#�ma�l�V]
ah�|ɪ����<c&{޻ l�M���DX� !��������(�1����lSH� ��ǂf�$IA�So�ǻ�9o����0�%�c����>@O��.�Z/�ߘ~�x�-���R*����'}}JQ�E�?�S>h�F5|5�#�<<�4)c����\� ��|�9�!8��Ⱥ_\��4��Jj=P���\�c�)��&���:UT���V�xΣ�F����ጌ
ǐ)��ܠȪq�W�H�F��YF�N����sx�)�%�6��v@,�9�p�x���Բ�4Х���}Ws���I�R:t��"��Ɓ�#۸�[{�,���v�K���a��}s��E�Њ��.N���9�b��;\_I��M{�j�J��y�ڵѿTUqrc�_B�As�'�(�b�*	rd5�gF�����EE&wZ�'oĚM[U���O����xȇ][���	[Hs���{T���}�%�&:U�}D���u�Ŷ����G1�dd#�{L#R�>�e~C��C���+�		�i�䩆&*���{o��)N�N����I36ԎY#v��K�8���p;o�ڣ��]"*��������˭��k`��&�I�ے���+ݗU3��#Cw`Ȱ��Qr{��w�52{�[q�4��x���]��q�HE���m���Ϟ��w>YE��9�AH	@��E�	�)ߢ�.~��m�-��\Z͡u�\�oa+&*䏂U�Z{ϥ2��h`�bް$fv<{�ٛ�����n<ؼ8k�jTV~�M�h��q{t}�}DYe>ܻ�k�0������SH	+�O`7��8;i zU����	|\�
IbK2��9���a�$޴��n��8��Ŷ��V��"B�$D�H6���l��8+�-b8 �lZ����4����`$«4>"yӿ=S�"
r�1�^F�O;MD ޞ6�be��1[3]���ڠe��N=nX�h����z�-l�!Ʀ�5+=!���7�M{��#�ų��zDb�2���ݕ�U`�wcʕ*�G���ţ\Sg�F��R���9e�:�ԠYA���-=b���(B�r�H��Gڃ��7��9kDkg�:q�eJL�s6E@�s��6����v��Hg��l���Q`�A�>�w1x|r��am�������@+t�]ٻ�zb�K���s�G��|�71�8%c[p�ۏH�P[��C'�2�QX��YI�V)^�u�]���b�ϵ9zΌX:&'f2O�����K�ᐏGh�q�ib A�E$�p(��>ᇠBY��D���*�n�^.��D�<nb����0n���3�I�2\�g�����-E\d�(�\R�
�t{'{W&��SnԌ�搤��"\'�&t�����e}�ٖ(�����J���J�!�|����z���-�i]1*����J�~ƴ�6�������m��]�O\F�/��O�V��e�kȿD%ql�D�-��jbQ��%yZt�G�#�l��f�Y���H#�SA�
g��(f�Bx�:[Ǚ\��\����b�A|�̝+��Pi��N�<pBm�K���8�y�e�^v&$�O�Nm��f/[��3�|軔�
��+𓉊��S�!ft���t���<�׌�(�l�������E�	���敉�V�V8:�[��pk�ø�8g=��W��3ŝ�s͂EJ*���� ��t�2�Z�:��G)lÎ�'*[^�	�:S	/�\��>t%C,?%�w���&��'�hdP��d�2�0�"ID�賴Ɉm��3t	�Hצs���J���3�J�x��DF8l�%�� �	��t*6�%��o��)���K�����\��r@+��!w/|B�"�(�6LAU�����;����;���r���:����[g�������Q����]���k�ȫ���k떅���k��\� � ؿ�Pz@�F���?O��*׭���͂el����hK�o�%�_=�p֬č���] ��K��b��� b[�/Q�(&p>U�G�_,r11Ѳ���:WBD���z�S�u�2s��T��@��%�[�*�J��6�� �	����e�C�D5DT��fW��<Ǉ�ݰ��:X���+j�6<PG���Ay:S6�M�$�3��O�{��Wi�^w�"}�޲�:n���2"K��\��+�+�̩4��z�E�7INA��dяa{ cR� c���Dq� O��I���8�7��k���k?�=!�oq]KGa�������xq�s=}`�$F�r�c^�Nj��PZ|l�fϭ�����`(��-<�7d�Q&��<พ���:�NTݓ�Ѷ�7����o�&���)�����H���f���֒)r5���p;gn�&�=�y2+Z!O���#�6�	t9�".�+A
?��8F�)+���waQe�$<�E�}Pd������
�V)�Y7R��$.a��ر��D½~'�4�f���|��C8 lX�5�Ӏ>|�>�6�3�>��t&K��vT��>�j{�rO)�<�&嶚�Q��]	�)~x����o�8BMuIþ�.��9��ͯ�l��+��ը�ES���EE�:�̠�k�ZS�4��.�nR�B�A.@���;�kH��n�A������u�E�`}��k���%�SO3ۿ�+0�Fp�b0�$��H��m�6NI��4�Đy��w�X*��i�|F^a�[Б��Ģ�{Fk7�L�!���fJ�V�'U�v[!-u�.����UZ���t�X"�(����⪠��E���v.=�}� kHE��o�[|p�Д+��$om��:��B�}��ؚ�e�AB(����K�+_oTb�C,�o4Y[$�@����{-j�9�$������ 9����''�n#���J���k�>ii?��*+�]%��/��C��\���\���ڸ�}4��up�x1�述e�Z��z-�4�Ű�=)���]�5M�冓?�d�^Ѩ�������!�x.��j�=�S|�����f¼�A�S>�f#����$n�]!�vz�����P9���t�&٬f����zђ��D;e�NX���M0�Z��X @5���3<���vIa:��M�tnZ�⬜╲��$�����h�C;F��C(����(�zsO�ٍ��
�*^�� 1*�4�#�Q�~�b�߁����l�i�'��/��D������w|���W~�Z���e-H�Oɕ7�q�;�9J���"�q:Ĭ��t��yM���c�:�Qk�)�K]ɑ�r ��$�����~zU�7n{�t��_����&­N�]YBI����@J�����W.,گ�ۙ��%����&��[��
��N��|AY�\��2ٟx��D����d����xS�:'u6	��6k1GMR��mk�>�4|	ؕ�$��|�`�M5�ݞ�"s���R�v�3��1P�u6�~��ٻ���-�z��c%ZIw�#�ڳ�,��8��.n#��:�M�z;;���������zC�^�_D��呾-�-�ܔ5��@��]�͋A�j͎��B���!W-2>W7o��Z�����g�^��X���`��Z���ϫ�
mh	7C��x�vgg���/���*��Pt��ݰ��#�\���K���+<�{S)z�X��r��������T��#�쉣�~���qW/j��V���(�0b�������bv'�ڿ�z�;=|Ņ!r$����a�Z��]�]k��%���@�K�
%HQ���j�W� �	��eo���eC�D�w���7<�nsgع7�脐`AJ|���~BB�E��8	%�*�k�qv��6ډ�c���A;��Or�hU�Z�d�"e�r��y\ܓ���KE��?����rّQc��W}W��U���ڒ�Z^�����"o�+'�j+$¶෗��tF�X_�;AA�ޮ%�W�|���n��a+d�r�I.�_C&&��!��Wi�W�l;� %�/O{��l	���鐳����y�?�5H�,޴(W����r@�)H�ؖpg��c)	�0���jKey�Y��4Yt~	�Q�&�3vǟŪ}��B_�At �`9f�v.��ʹ��}�*�?��u�N#���gI{&#��.���G v��l��Zݺ�#	�����2K&Pb�aɡ�ӻ��CJOE-�VV�g ����
)��m���ͤ�1�5�/�>��Зd�"Q-&"vMp�I��?A��9�VC�Ҍ���StG@}�:���Dq1դ3�3EI;
�`I?+���`A�3޷
�}�z�1-hu��O1=:�3��	��=��)@"\��/^���*V�*fj��ihb&�R]bK,W�pNS������(=q�_�w�4�#J�tk;���'3�����9+�l��;�o_���pe1'u��RRb3�{�E�lǖ����P������6&���ض)�r#��峀(x$!��j� A���JwR`8��6_a_a�������4`2�Ŀ���f=��vc�G��YY��s�w�b�}b՟�<�!��V �����1̵M_R�uI�}|fs��Q������h!��o�<ɍ���)�(B���5"A~\���^&��c����$7�A(�^�WC<c�F���,�5�<�	ѹ�-�!˺-��Þ���x�R�����3��ޅ���r��xVa�|���$��,�yc��s	�B iJ�u��������u��&�ɗ���m�B��2��b�fp�X�Tt(]:�S�r�i=��c��~n��9݌7ҷA��1`i��`=~Y�)>�4|�h���iI�zr��v�>�,g\&���#��	�m9���?V��b	���L)D���G��꟮��J3�Fǁ�#� ��1đ�@�"��˨�Xz�o������M�`�V�AM�{�7��ʪ�S�'��o"
J����(x�����6~�'��\���� Lv[4T���~��;S��]��]��#�	������sрBf�I�
z��U�%��Ho�p��ݫ)>�{ߝ!���E?�:}�>���3E,�1P�V+�e-�m��D���[hN����2����^"'����A�$�~CW���϶�M�/� �tP��9�(�NL��A���d7��4���V�chZ&&XC���8`I���{��i��} �Ybx�yG�����f���d�^$��?���R@�P(��>8����߻2V�~6�gb݆��}t4�>|�C��f6���S���e�v �(nmLbpe>ґ!�]$#�E��,\��_rw��0�v��E���w#U�����7U�,l�v �����J��Zj�^����4 ��3�ɇ��-���.
`W,܁L����׫q��7�_����X�4��PL�<�0���Xym��}l�I�hkM�I���1�<lmN�E-���`}���M��~ �yCi>���CD���l;+VD���)Ĵ�Jj�L�>��Z�y����8B����`�,6 �Њ�=F;枋Nw���"MU�"�&�����iז��Bu޶W8����E})��tݵ%ح"jSa�-v��vg<4�*���^0�@o���^d
�4ք�=�+r�jrg��IFn���ъwҥ��r�P�Ϛ��g["�,dh@W��9�oA�,ӧ/��~x�$�{��ʰD~W�&�3�N�B���V�!�y�P0��s�n�?������?M�r�}Xt �U]����~G���}�S��]%�Z�j�it_��-į�����9��s��3�B�Cg^�(���[J���:v��� ������ڍɟ�?�τ:�k�@b<�_�ު
v
�N�]W<G���9����7���D�G��-�[s)Z0��J!P���·�E������w0�x�E��T��*����e���& 2Rӈf�R���v�fܭ0Y�ҩL��B����F4�)XS�ڍ��S��v�4����
�7��7J*����^���1���Tԧ[�-L��F.O��C��E}I���y_��M�<` �s�܊$n�UBu#U�i��]��%K�&���[sl�et�I,۽)-�_�g���Te�嗒�j���o'R�H�a�;J�*ݒD��1'Ũ.E��b�W1�1�P!��oij�����*E]��j�ݰ���}&H/y%{��CU���S��(;DA��01s��d�z �)�ܧ���<����$��_u���V�%{�X��L����Q:85�s�H��)�7%C��AU�o�$˶D�c�4tg�B�s�X�Ӓ��k�m���G������l�V��-�RwW�/���j�8���z�h�4hמ%�Ky�&���g�g��K��)�W�!��}=[��m*rIj��� |���D��|!)uK(���!����<��0%�k@;A<6~~��#28��P4,!΅����G��zz�I�h�x���'�D7T;K�
���ɒ�*SI�(�X�b�ۏ����3��!&��(�I��؜g���Tx_fFS%~�"�?�`�ƌgY��K>o��4�[�!C��L/x4��^��_zE>j����D �/̣ ��|��ʺ��o����:��[�j(unNA�i0�9��h=z((tK���N`k~�H/g�H���M�L�}`���eDC�2
������^�ai_�%C��3��Ƨg�4^9�|��@?z�*��]�P/�R���_��e/� Ȇ�'�r6�������^�MgK	`�{���z##{��
�ӄ-��7��J\�ͬ����:�W�F�h�!iseU����N�4����nNY)��E���eϭ�΂x��)���\���J�g���%V�e� �m��M��(�Q�7����bS\*QׁN��y�j\��bJ��|�<~�1+�>�+���:��w3D�/o�>%��f��nl���Mw��q (�Fy��S��Z���� �r���&|c�wp�"ׄ����rP>���U��Mq��~ē�݌�	qro�vf�,���d�*iAV�U�{|�w�U�#��kP�T$H
��1��}0_[O���LcFF/����H3uh��?=8R^m��Xo�Y~�	F3
!-5���F"*��9�f�;c}��œP��S:�%�w�����5�^��)Y��	R�ͣ�Q�gI˚���Y�#�#Cr�X�}Q �+;x�ݞW�yyv�A����rA�t�޲<G�	�u��)C!O�oj��߻|L�髦��\�E Z��_�û�EZ\:�#8<A-�u,?r��v"�S|V�ە�D��&��Č�
#�F?��.݄������knkr�Xd�.�"�z~���ʞrH��S-�T�����nv)��E�8���q�$�b,�,X�=K��_á��6p��s�!ܴ�B��n��s�l�l�D"
Ɉ��K��,��f����h����d���EQ&��L/bC4�W���nz��z���I��=l�m�NZ�@�RQ]� ��X]+�`&G�ZΕ��dBH�Ò�|8���Z�v!�,1:���4�� �ͼt�����7j�#_yJ]wC�VZ�z���֙�vh�5TO�� ����ݨ}j�pآ�S�
�AC����,}��iݘ
�7qP�*���õn���SM�&�e�Z��Q�Iȣ��[�e$.�<�;V\1$���5�ĉrj1`H�&m`�*�Ev4��т�3o8��O$���=Pu�kf���1!�[���gVi��s_�Ft��"��K��\� c��ɰ���w{p��N8e��ZM�'*Ϭ� e�_<��4z*�����1�k�<��^,��o�y/�w�8������Ա�SyC2O���LypP��o�֫��D�JB�c���=e���E�*e��"'�,F�H˫a<mV�h��%�3�Z��"dtOe��Tŷ�F)�cSI&L����kx�yj��n��$*o<8\-'r�g��j���̧EU<�Mʡ�R�nU���ұ�n��p�W�ʻ���Ӭ9;z@�����P2`��^^Z�� �%�-�&=�4^!P�-r�pM��\�����#Ⱥ�S�ձ���F�&g�i���N����&����XMNp �0B������n,ս��C���O��8�(��
S@����L<(8�l��3X��V��O7遆�刭���7,!��!���Lw�#�_�!�Q��[^����j�&��!c��C�M������x��&[���9�ǒ���k@���|�LHm���'w��wa����괍]�T�GuS&`H�Q\���щ#�Ooe��S Oɩh��={��!�}��V|Zp��$�i�KS�iZ��=W�%�cY�?-�
 �p-�!IhX�u$��Qo�{�(��W	Nf8���A\Nc����p�v�Z�}װޗF�Q�|�������!zӨ��r�9=K ��艊�<�G�]��N�&���!�����OeG�-�MK�������`l�)����X0J��0��sK~ǒ����&�]�4�S=ǅnҦ�a��>�=�gL�:`;5�3����g`!N�`>d^n��3��6u�����)Q����VZ��=�2O���$��'񞓝�f�V;y�RB""�����!W��Ϛ���x��#�Q�8�rG7[���#�C���DI� �2�ZbwE��}��8�r�l�vB1I�?���>Ȉi>RP8�~K/*~�C�P۞e����]��7�p�	H�����]�˭s�d	�+H^�M��ª��"�
�>v^��.N���:��w?�Q�0�G��W=L>�szs�b��}�|^��M�-��!�)L|K�?+�2௓[R�B�E��Ժ��/��prIk8za|M��2=�1�Ɩ����>�&@.0a$�����j�u!��F�k$cF�
��⣿vi��f�gF�����#�Ӏ�	���������hA�..���
�'Fy���B�g"���Ջ�s��ڒ����h�w�$�e���8�P:�4�E�w��K�Qdm�:���"�q�B��3��{�$;"��-�W���/���Jt*��z~/
|�mx���	��Ō{4����*Y�|w���X9(1����Vh�b�|�:F`"a���<��9��$`@��X���T�f�Z<��ܝLTt�d������{Ш�)"� fʅ�"1��q�&���=o3�}5�r9vW_���xHaHT��ʏ|x:�;u+�]J�fk�`ϜE����eB���IS�г`���T�o�ȯ���I6_������ۚ�;��(��'�����t=�e�ui����Z�������+����1��Ng���f�ƺ&�u��~�\{S\��n��:4���f����+���>K�A������P+��a��;���5�oq�範ͧ3��8���u�^?-4/�9����(�4���;0����Y��2r��Jy2�@�Ҋ�R����M�A�dD��JM\�w'��:��ss	�����/�Uz�KQE�3m�~��0ad0%A@A)�^Lf��g��'6������)����h�O���V'�l�PwM	�
A���k
S V���D���R���(Ino,������.�\ͽ�Ňh#��ޯ������.���6�.�<�����`vRs��X^<�A�HK��4�We	��:R�)���V�/� eә�w�2(��
�tR��>/Ja����D�ҞΈF�b��V]\0``~�D�t�|ctL��EfB[.7�הP���X�������l�Ef�.��"o"�]�-��{��l���^��f�b��l�V�̒��i����t���$���G��ǚ�T��o*"��5a�JN��>Um�.%�d^��I��A�59��'��C�����ǘ�2�v���4��՛�<E~܋��?�FPN�!`�#�2�d$2�Q�&4�����<E��Ded�b./�\��^�/L�R^w	�(����%������r�o�ת(�[�S�&w׾X5��A6��J^ƲMc7ע�mWs�ue�1a��u�Ώ�
]�\HzR�����qj�P�]�үD#W0xk�)����U�ZL��l��5[-��.������fo��/���'z�7��b}Y�nC'��'}��ì�=��>�K];��x>	�dx<7�[o�X���������>{��������ز=q�Ł�(�8�;�Cٙ�{G4��s�r���g�tģ.�����7���Ui�g���pV���} ��v]�ņ.���o�ԜJD}U��j�8��q2Nm���]�ZiY	��rYe�Q[�y\~'Ė�߫�Iݡ��6��ɂ~��t�:PE�<�)��m5zK����7����q�����4�������[Qg(i�K��_�9�A��hޕ�$B(>��.�J6�)�}c`mT
,��	P,z���`�-n��1OE�
���\e7;[O24��-9Ø����95�9�V퍣̓G�Oq^�F������/��0*K2RCB�����@	�a�)�G#=lЗ��5b�`'�-�N���R�A�P�9��F'����eͤk��)s� ���ɋ��G<YeLv3�f(��>TpO��@��Z��T�e��:��:�D}2t���R��TH�$���\^G��������P����m�mmY����x�fy��#����Q����?Q����
AK�P?��=7�u��Rqe�y19\��BɴA�x]�#iR�������:�{��9vC����'f�;�"窌��"�j�V����P �#~�._9�� W5�6x��jr�JV�h���O(ԃĖ���95l�x��I'�VX'P�RT�F�p�C�����M����#(Ѻ<���a���x����'fT�`Ѭ�B�Y��3�����wm��V}s���෨�=��̸��t=h4�k1�<@�n3��0��*�6Rq���{_�%	��+$����qSF�\ɠ@xЮ]��F��̯��Bel�(���𺯪 1�"9�#��
b�!��͔M� �74��K���@�j[�7H�,��n`�;��<��Q��T��t��anً�68�54�����bE���Ѻ�h�yG{����.7Yn�Hn�a�qfP��g=���$h`��3�p�1\
��O�Q�9y� �'i+ "P�a��,P]�g����u~Z9'��֠ᜒ�R��
�a�xO�ns�<�@o��(\�s1Jڵ�Z���c���
>��'�[A5;b���/#l6^hѽ��W��|����@"tN٫��o�+��&Dڡ~�!=H)�s���|6�}Bm�5E�|jCqY��F���_����Ryi��@RJq�V��6\�]CA#��K
�m�&��k�qG��w��4׆-up�D���߱4�I�P^����Eρ�WmG�	r|T^�ŃO�Q#�=�2X�	?���<I�*=�p���:2���V��:Q	��"�C��Լ4 L�Gf,���s��ƒ�/�$�/��g��6@��`+	���D�AkȜ�(���������Q��{������2��f�;���1��H�Q�/�{��w���x����LR�{w��`���@B>_�q�q����?F�a�%@$�9�IC�\4^��.�W2����FJC2C;C����ʚS�n=>2Ҍ�&��鿂�tH	o��;2�p�Yu��H�-�`�k˺��)��u�|l�9�m�_��}�'}�Ά�1ש����O��{} �r�E�����r���(�Z����(���!�_�{� ���t�����/y��+�|
�s�����?Fw�vZ
�N�����	�%�"�Vφ�{��GЌ �L��
�xY��X��1�֝��0\�
@����X4��Bï�gX1�!�8`�}�i;W75I��Ak��E�(Ad>�Pa����Chǎ*�/��`�H	T�{�;��������f�����r��'\�Å.�'w� *�8]�t�y���LD��$��'b��!|�0S�0�x��_�N��v�^nN�ʴ��������"�8�4/�����SG��8�{{]jH�ѝ���>(D��_?��_���b}�������h�+L�o��ʲe��N,���:,�@h�&�]���^�]n�k����� ܅�\���΂�I���_�t�M`)��k���IU�=4m�	�&�8h4!:��4Im_�����DC����&����6u��HH"���N����+,;�`0�Z��X�t��h�Pcp,��Td?�[>�t��f��,�Ee뀗�e���>ߓ>.WQC,�F/���Z`��Lb�$�ZV�L�Y�Y�����ʌ;��걥N�,�0�y� q���L~5so�]j���V���X|��u_t�fm�D�&���kE���KW��-�~���\H�tA 1)Z�v�R��Ч��a	�xL�Z"6���3�E����Cs+c�q{H��@a	��A�ZI.UR�Q�[�(��v��dm��㒏�b�Fr�b/�5��6���t �:FlZ}�4���+~������ړE��\�� �D�ko��6o�KM܁ϵo0��r
Q����a�k�?��9%�!����`�/js��VSe+���F�^���K�p�#��!���N����ЩUV���1 v6l��\ Z>�x&��������Ў�w
�1��Ɛ���q)5��V>���<l����&� �!Z���M�q�\6����|څ��ma���o�{#��Uȧd���R	��p��YX2�`6���y��+�S,���O���ʐ�*�S�:D�)L]�����_#�a�G������9�3����O�Ʊ���n)V���Z
^���X��M��I9�Ha�{���v�[�ߓe��8�Lk���������%���؎W�0�E�o�4��R~Sm����F�����ܓĳ�\O�=-��NMkh�@�M��ɂ7���~����-'�5"��1?��lfY�٧Z�����@  �XGjҘ�����X(De��q��3o9���.X� ��4=�V�ɝ��<>�Bn��Wg{�O0Y�B���=l@j7�^7�V��1�^5dL��ǽY�Q��e)��Z��040O\�O�M�?�Y�#�����U�)r*��d��u����H��1�uY�Zr0�zW�Zm�kqj�~�|h~��"q0� խ�3%!��,��������&�?�s��� 9}��������9^�$pL8\��,ݙ���4����~C������8/+�Ҧ�-�D�ì�.��喰 �1� �PJ�\	aM�̝�^��ʎ�ɐ���D��F����S�I6�,Y�Y��kX���\��(��NY�xttr�խ��Ñ�o��DIi�Q���[G���
Sr_��h^����ԅ�Jc��ϐM�.`���w���w䛺�4X���FdpXS�Hx.�`��7nZH  �4{O�O��^/��1��k@}��%h>k^����]֝۽��i梊�WVyQX�Q,�}ɇ�/��c��M�{�w��:�Lr�~'�,� 3*$^��nz+5�����N���)E�g��"�Xg�0KV�4�_�bǛ����l���۸F=<��I��k�a��Ҩ�9�t��08����-ғh�#�ؑ�z\��,rjr�c���&��eE]�:RQ�3�A75�I�-a�������~�G9��g~��Vo���8����p!�&s��s7}�>�T='��d	 �_��3�ck��;3Ǿ�(��"�� �#��з�f�2��e�j5%�l�i�a���w�bHzM��@�.�]Eo�}��^��)	�0A�~'
:�nkц�͡��Фsͽ�?������Rs+��U�o�O��|���22燋�Ȧg���UTCذu�u��ÈGs(qV��Mb���a_��&6��]����ò�Bs�͈�"�9|m5<�tS�(2r�����f��f�h��N�=g^���¢F�3���1[�v u�1)B	��) 0�u�� ;sP�b��M�=��(%g+
oc���.M-��U�e=RE8W���v���?̴*��􏓸P:��F	T�[��s$���ߠ���U5@�^j�X.�Nؤ�nT�ǘ$������?�4��k9���0�ك!*'�0�`�aMӚ�nM�$���&~T��n��J/�̪j�tҋ~�I�A0T!�}u'Q&��ƃ'�G[��e|q�������8�Xx�� �
I�'<�f[�5�I�_�d~���`��X�&�?	V
e�%K���Ra�Bݢ_�N)II!:�k�FX�z3H��"8�dN�w�K!���M �a)�UztN�s:afD}=.�"�C�����I����*L�AOVK�(��}sm��hf_	lq�v�n�>5�Z�Gn��|	�V�`_�R�/y'�����b1n�33��ޱTR,��"�^E�u�b+�!�v����v�����L2�|��#�|��	�گ��֑�I=,ؠ2M�Pć+���7k}Z�ǡj8/[�����c���h�sv�=�6���/�O5�
ʜ[��l�N^��#Vv3M�K�z�kK}�bg�$b�a�u��ل�cE;�)�������6Ɛ\�;/k�2�e�����!Q��C'è��v+����bE�5��<۞�E�����TмϪ����/r���\��V�,_�Y�1�=�$�ޑM��؀=�%��#T>ݚ <˶S0B�R6����kH�+�)��pnܺ��c�@(�8���2��^v�T&,�K�J�����@���#�eK���L�H�=�m7��_7����X*��������U�����'�����'f�>|�8�J�V���9ˢ+�^a1B��,V�0�7*���&,4����0Ş�n����ĉf+�y�#	��Q)����px�+œ#�]���OaHU��-��7���L�����{b����&D�u݉��]6�|R��%�(���b�[�rC�\Ӛ����o��a���~�#�+0�-��$0�͜�oLl�[��/d̉��
ը$�� ~KR��a>�Ԕ�tx|�рW[�_Q��oKg�J�Lp�^��x{g�?V�|�QR�W���9N�}����v�:��9�8�x�y`.�4�q��%��k�*B�߭
��ϫ��G ����z:�U�!pe8a8n��:j~��?'f�ӷ���������Cf��K7�h�sp�>뷦Zr��.�CW$ɮ�0�i%�9'�J���Fy�D����U��K���m����緎�h�~vذqi�A���TrL�iĪ�^���l�W@{eѳ�L���r�TD�AK��h�����#lZ�}V���cDVHQHz6�ӈ���5��t7[T�\��t���Z�R �1�֎��F�хu?��r�B9ē���˸n�u�#������Ӈ#�V�17ǷJ�3�{	#��5M�6p�AK�y]E���o+�W�HĈF��GT��<��yi���(�����.#�QK�S���-��YLV�$�|��	����4>��""�ĲT8M���S���ϯ4Y+6��&c�`�s�R��嵗��'�t S<��˲��
=�p^U� ���hFj��W�{�������:T��/�1|�S����D_�	s�d=Ū�*��ī�p����q$5֠r.�ת���l
�D�-�:Ā�Ie?�M��$�D�*Sc�ܰ�{-~@���,�[��M���!d��OQ��:��dXC��f*�Igc��`v���\Z�^oU�ם��c���ӳ���RT��eε�Z���Jc#%w�U݂�Z���hgT�e��}e}.�u�馠D3����}�"�f�XF�f�
A�I#��o\m�^��q�G��A����-��#�7��Lw��8��du�G��Y�PA3R�	@X��C���9�"�]'6��Cr�q����	�؍�jY�sV��3���}/BE}��ĠI��!��,۬	�ңt�!,@J���1� �-J�v��R�j���\ �����CmV�A���6�N�Lm�\�\��)�/m}�Ǣ>GsJ���:��¯��,�Jie�BC��gu����Wuc��%��s�VB*}���u��EOlĕ����[_����qv�<����Ű���K���o
hV�}0���7�$l����u�8��5om�&��O�J^w	�=(�RH��M�b���q�� �)�h�`V�O��igZ^h��=A���0�)�����������no��3G�*z��-��\\�y�pb�$�@���	���v2=�K5�o�0U;X��7�!ʣ�=��X�ĭ�=�ޜa.~�ٕ/�	K�Ayi��+@�->Bw��,,\�psD�*�P��'@)$̘]�~�f
n�{c�Wg�V���"�GڎHɐZ*�ClO:4�'j��]9�O�aF�!���� M	�Q���89�v3�*��R�Є�a/�}I�_MAE�2���I�5����!�(N$�����< (T=��� ��~9�XK1�7�/�T� fʺLщ�^�>Ո�����u����x<C˩������{:���my�~;���fY
. D��"w�Q����7���wl�!c��F�yJ��%q�	"9�/��2rC���E� �-�<�+u�sd�����t������j,,�Q놳����#�?���t.g��	�NͫV5~9��_��e=�F!ۧ��
�r8��(3%6F�G��D�XpXtL��
��� bAN#Ə��\�TV�'��z�J��f'ֺ�ѐ����͑+=p�$�d���{G�b �ȵ����}s�9h��f�(��A� ��V?�c2���3�{�[p�3I�Y_�`�V�LUTd�N��+�����w��L�\�ׂ3�>�ib<���d돨�wFw�	�2z8��ܜ��T����[��t���.ጉ@{i���]4�'�P����,=*��L����D��$:�-���њo�Av[_��}T3�o&@}�?�T�Y�M�0q�Ehp+W�/��ݝ�M�� �%�+E�h�����e�Q���W�rE�p���a��W���غo��:���ЯQ����f(�V�U���B0�!�Q�H��eX	u�NK~����H?>��k1�\$\�>�T���<�\�!�%���0c'���b�W\�O�H�7�h� ;�����Wp?|����T�b��U�D����}�xi������}O�|m3S�߱�W�p�) %.���ˈ�b�*�"��gg���M�� �|�7-� }=lp�����]�3��G�
~�#���?�M�	g��U�r	�~G[#��?¢J�9�v��n��K����fU��g�N�m�fA�}���Iƈ�P7��P`��fT���~n��V������0�W��TAQ�KCD�0�~��"9����1��Ds-� �k�!���&�W��C\��U�����1�����|$��?I�x貧�9}���g���z;�gY�����@Qz�!��ؔ8��q�X���3N�]d/�y������[�\}5[矌�ѡ�#�9U����iÎg�" �F���5/4�:̒4��m��:� q�r8O]
b[!$]��%�)�d+�4�-DZ���@gZ%C�Mt�����_� �ƶ��f�(]�%+A�j�\=����0vs�-I��r#>����B������Vڛu`��*�H����6m�@F�%�k��i�nO�����R�m���t�p�ȕW�ba�)�K������x�n���XSį����Ҿ�d��y���K)��`���~J���M��4�h칊S�C��������bf�.�y�N1Yo1��C5H�g#�W�8�Pvh��$o>�2[z���>���q1�6:�2��|)�� ]��׃O�Uv���)�%y�R��R\�>�'ݲQS݉ˈ���)<Ğ�cK⿿�6U�Fj��jJ0��vTV��<ȸp��j���!i��oE��^�@��ˑx�ּ��L�2ֶSD�sCN���(E�O�'�STf8H|����*�(02��:�5��@��pO�9�X�V�D�'���M`:&��bg��P�u��ŧ�b<Qǭ�f�)%(~6#�X���
��,�������[�!D�@��28�(��år1�ST�/UϿ�NT���b-�#������Æ�A'�s?��-����MȞ�sK�*�p�6��0�
N/����P���-� A�����HI2w�r�G����~Zg�#e���M,�4����0�h�����Ɣ��'���'L+�rLd�U��e���@l�-i].t�4��'��0t��1���!AgIqN~�w��?g	��o���Ь �a6�y�=��*�8`:M��Um)~��sޛ!�c�E���+���o�4��Q��[��R	�0HX���ShӌB�8��	���D��m�O=j>��*���i8�5��0��խk�#vǂmQ�(F�9
��$(�G��}�� ��%��6]Y�\�����Bv	�[:m���X�K�kl�H�]�<C�̈V�M�t�X�"���x �$����SCT���SR��wu�}�LW����5d{*�n�1�?�񿵭a�4�̺�g:�X�&�-V�[�,p���6B)x�hv3�^�
�+,�и�.��nA�5cF�"�ʭ˰#�J"�?��/��4�1ݚ��;8b��Y2��
��x3_N�� ��:�Gsx5�y�����:�����(� ��Wu�FO���|'a��k�W�@G�<G��xo�o껂��C�=$��[C���� ��	��dj��ͯ��ğ4��}Sx�g��H�(�h�x�_ K,�M&Su,߁L��@��@�X�@�~>�I��D�G0�0���E�i����){a��ȩ󑱃Z|�&Wv��Y
�X1r��4A<C��V���bw�@�q�f�T�\�q�U�*AJ�qwi�5�x��KuW�,�O֫�0M�����̙�_Q���6Q1T�mT|��}V8	$���SQ���[VQF���]P���\�[-V�����^���������k���}Y��Pk m;�3�3�S0[�� �BX��TG:	�H���,�	�mϲ\>����~��
�d�4�ꈄ�2,�;�����4�ǆ���O�[�#�)T�#��'��Ԗ�7=�����[�s ����a�tod�A��qt��>a��`��|vN�Б�	��B�ITl�0��I/
�{�s�3F�F�|����]�J�if��[���;��U��l���q����Lb~��ь!�n���~�Z	W6��^$�Y�?��e9!��� �d��q���2ȱVd |�\��������(]�Q�]�J��h 3�����Udu���;�ee��N�|̭ĸ����;~Z�*�:��F������	%��B�*�,/�V�:�#9�W�"�+���|�+�=�B�d-����D���uU3�H�55����J��u����d�����a%��T*'�z�99�;���֭]� mP�e�5i>F����y�P�e}�G����Lh�{��4oO��= ;gO��@�<��U���Uz;9I�8K�P�aF�1󝽺��(B�(�1�qI�-R��i4x��E?p�M�a=�����W�ۖ�k���Pﴎ�,�g������w��,�8 0s����؟�ٺ|@d`�N���~f�m�a/4�I�{�c�F�^#&��w�;�.L�)ɑ�=�-Qg�����0e�rjl������K��{��\��U�SYdQ`���-�|�sN3�Ŀ���0Ğ�
��(�m�3�?�N�F�fr���pR��$,@��$]�b��io\�R2���L�C�d dl|�>�l��0ڛZ�˕�b�i0�$���{u�~�^�~/�=(�����:�}DZ�q����}�O^.�Z<�.��UmT���7����Ej���u��W��XRFv�� 7����~A�=m����<S
��mq �&����q)>-쎜G�'�`�F�;T��AaJ���%������:�;�(^x�*;��3�k�R���$#�B^A���@��R���U楠rx�9f#rc�ʃZ���Eۼi��f�[\��=W�BY�.�1���W�L�Yv��\�x)��O�:�BePVA|��!��ǰ7(2�clI�_��b�K��^	\�w^��1S������0�#�\R��P7*ܬi�~�Re빏,1ւ@В��3���d�,sA��~n����e3"昫v�5w�n�!��~S�#��/��l����+qٵ�s�@��U�YM÷�F͍_�K�6�`-�U��\������,��]&��,0ή���g\,����?��A)�|�+?'ajF׫�,b���(䪊1�DR���ۀϱ��~�������r̦��h8��1S®fBL$�	���F�C���WBF�&<� ����I��\4
�p�JSV�^�@6kx?tkw�׾V��7��N��;~(-����=�f�>�lw{]�����ޗ����b�\��'āv�>����.�(�H2�Y���L�SX����N�W��KQ�f�L\0���n3� ��h*%��e�X��v��̼R)���@���YvARgF��-�0� v����ֆr���\��2P|��ˇ��8yX���*�+��}f[n��Q���t��(���A�˙-��iZ�AҸHپɾ���9E�L�T�{��D �V�%Qp�:s���:�40e�ծrY&�<���l�ڀ�deYIꍋS�hh�(2�ڀtvr��Kjt)�O�@�̄�О������5v��eE��nw��*�q����⻥��|�}���k����nq�)߿{U����W�	����,T���[Ťr@'�&��%�k���h���5���RB?=ݵM׆��LE�s��s���U�zK�O�%����}&�u������#�)T�>�Yt<`w�п���|q��kߍ���a:i��\r%0�EG\���	�f���jq�����݁�Oz���?}YPL��.��Q�qj�W�}�|,�\� R�,��l�2�I0�|gή�Lb��չ���b��fY��z�D�����S�+�V�>2�
R9�+�"��F9"",)��$������;%������pr����>���i^��t�ȵ\W����N'�L	N�����
^lX���!6+���+pA賌���g;�����7��#y��)QL~(�����H�I�Zi�s�L�X��cM9�1wg��[�*���Y�&��yAN�op�� Lfſw��zN���<6X�0���,�6.���8\e��642L�k�Ii�
��[��>�@�G���[b^�%<o�3=�0c�Tq��V0��ky=�Q��f�JW�i����V��Ĩ� ��nl��{�F��0	[�)"��[�6N;>ҧP�|4)Q������i{#��[Ȭ�tm�vK�:6��� �Ɠ���/��r`7�x�F&F��l>��@���As-��;�xI�i|F8��<[��!�r�K9�9�ƅ����؜���
�����2�_�����n<O��7���]�mWmz��;�B��Z�zD��8#�M�H�i��������ۡZ+l#?�$�]�h��y��[D�#7��H �7� РK��:����y
g��^�ڑK�xǛ?Z�6�O������I��r��
�ښY���t����4X�j��dp1���3\���TX��Q8�+����|V�/�ѳ��q��h������1c|���=������n���Z�������bΫۗ3n]���ji���q��r�f�n��s����o�n���m{�<�C��ˏ3��W��^����q(��P����j�\��n)���*�j6p���Ig����ܟ}]Iːy��˒�����8��EU�b����<��y"��kTPR�'%�@�B�t�0�/1A0<1ؤ3�o�s����c�@2O!JpOyL�3��i��-��l�u�Bt��h�tL[��fs�
�Ytzv˗�-HP<]a�Q�NR���Y��{���RIB�-;H��C
������o0ުN��f����~�?���:�ސe'�r�(錽ܶ����A�K�����ɯ�d��@D4^�\)��M rC�DNS��kdJ���PJ�p�X��r6"���^������� 2|m�Թ����]�����t��C� �?V
I�@yP���)f����*~;j*|7Pſ�ǽ��l�P!4�F{p-+6��s����L�R�W��CJ5:���A��W;^$~70?f�*�(����'b~�����J����Ĵ�ty��#]��ŰӅ��lZ�K�>���U�ӑB�z�"w���C���az�O���NM���Ue(Fkc��ǽr7���o[:`�AUN3���A_�����f�������|a�^�Uj�|=���ݬEW�	JZ�J�7B�DZ0$�f�H,&Q̡	��z�9��'?�sٔ�pt1���ڦ�}o�1F���"���z;*bL�0hl��8N�T1ƒ!p�+�H�"�R��~P���3k�y�#�<d����﷽��:��k�}�ˑ����ۗ���-"m�i���m~�C����s�9��&���T�o{�x�H�Zl&���p���W%�kF��,�W��%���<fJ�����6-����c�sC��Y5�Xٸ�:�� ')SO�7=[jK��}a�'b�gD�d�����Oow_���1�u
�!�,�d2�e�,��<����}'�3ZolN���\5�`��^�)���%�O�Sg�~?.��[^�������`ǉm�`:�L7��ݓ�M��bF�6
�#VW��C�nw٣`�Yȫ��U�^�V{+�:�x��8p�M�ڀ3k/bjԃ��l+�Д_� &�ȕw#�����e�Uڸ2�U�~RA����GW�6,d�����4�8#ؙ;iS	b	�hF��i��0'�]���Ss�Dt�?1�_f�5���?���&b�6%L7���v���<wb��.�k��]9؃��o�`�X��Z������$];��-�Gs�q�I������a�#�?)S��s�"\yE7�&Rm�U�H'��?'��'�Q)��2�9�7ʬ9�XQ�%/1�6'c6m|�\��Ur����b*��p�\���d �aw�:֥�q�H��v"	1I!)�(�O�`��w
8�^��0iP�o�4q�+	�rf�`�G�7qk�!�TNN2s^���O��=}v/W���J��D�S`���݈���E���|�i݄����~��dX�hl���7���� ��6<���@Ґ�w���;�;���������1�]5҅�k���2d��	:��{�ϊn��-�\G�͚�p$d���C~�L�d�9�*s�(t�~#�3�7����>�s�+�x�h�.�7^���p[�kE-g��릙7ǎ=?�U�e����޼����X��,u��s����{�������s�^,H��0]pҸY�ƄQK�n��p)yl��C-F�4nc��x�")7w���٤ː|������v��)dU(�tG��+D��H��Us]���#z���3�f�qF9k�'�'�ȅ�Ȗ��(�c9�xŖ!i�B�t�HWuH#O$>��k�e3	A�(���5�����6�Œ�]�@$� ���O0&Bf��i�\��n�Yף�y�{6����"�``�!���=�b���'8�y�fl��{,�}�W�<hwK|�?����'X�9,Ƃ�b��A���z�����0���,�f.7��S�����M�b�K>ub�ٚqW3�q�(��X�]�.��F0U:����1��� �5���K?�ʑ�1�f�ɕ>�L�I}��+�p��:B�Wd_��@@>#X�|�ſ���*����	��S�=�Z&[3�������َ)�"�~3p�=O�ъhu�iS�:ϳ>��s����[��^�cA|ΒU�GƗ�ْ��'%�Q}tTkZw��$;HQ~k�z�ms;���&�Z�>*�	�I�3
d??��ra=|eXs%�2Sb�C,6������.�aV*��N<�S��6X"F�T�k�R?��G\�A'��*\h�Y��"�CQ`�z��Z�^���������b�v}B�E"@f�3�D֌M���xK����3�9�o�e�1���䍺eYr`�o�~9�{#12�&��尲�Z�ȺI�v�a�~�QN���R^(D�F��"�r���FO���O����D,\�5�aMaki�p7=�b#B�*}�|]0�ҧx�6����"鵴��Ɲ5�
���+����E�ީ�͛uQ�~\��O��F�3b�&s�^��m2��y�!V�Vu�J�2:�Y΃<nU�[��ӏo�ja����$�����il� P�
����R5G؟��YR�!����R�Z��̀���DY6����`�-$�{�@��=���2ɇԍ6�P��O��V4���v��hsY�k5W�cW�#�o	#�Խ��V��ê�C�NSp�6��e�ﺠD{�����R_�i�+b	�bˢ`��>qqPJ7 ���qb���.������udf��� ��?h�V$��|AIeEdna˻�ą��-��6�0�%�a����&?���^�L
��q����5u�u[I%�T��^
�j^м�Wf �1��f�"��?򀎣����kr��}zeE5r�z:@ͽ��W������)w[3ep�fa֝�:ʏ�:�KX�Dizh�\_&B�.H-6Y
)�lXQ��{{kg1��j8
��W
��k��T��C��X%��T!��u�杮U�|���#fP׫��Gsa]�V�I+���\:(�@j릏��N3��d�0Q��=`�6%-�������������ׇ��.}�9q&Ի�
Ջ!���Ɇ�a�Ԅt&)sg��K��v��%��%�y�E��}
2�DǍ�ğ5��*7������n��q4�
d���-	+.�?�c��SC��F8�
<�O��ɑ6�V��Y�p�� G�[�4��
!�,���m���Wob�1ut�L��ё40D����7�d�41�I��9	$�I�ġa����Z}l� .J�@����l�n��X6��Yө�o}��C�%��q�G��_YPR�E�*'YުI.W� ܑqCy��4º��.���L+�u�����8�b�q]����z���"*�b8ᜄR9��i��;o�#w<7��E� ���/.$�po.�L��*"����S4�d8�̟m�I-oa�1�E��ɻn�d͂C�Y��q�GlOn�n&�R7/P��
 k4+�j��v�_������}*��Jl�|j�褂S�]��Y�}�Gr�<����	��cC����~e��?���Z�AAR
� 4�8���-�߯c���h+��3G���F�]DM�<ߐxa��K�{��JM�F6N��4��rrl�9��q���Km�bF� L� �#�b��
�-ə[A�>�Q�P�n`[��^���0��r�,�+��A��-��r�6���b	����}�f��x�a6r�6G?�����g�����Exr���kk��	���Si����f�0MA��uc�!����9�X��uk��"��_�ܠ�+�xv�\*��{�v&�6�XH��$��� -W��@���ͷ�@�����B
b����a܋�c�F�͛��F"�o����z���"� �X����<㵋�p�C�V�N�ľF:��Oⵯ�А�/���ć��Z;�~��gu�K�C�7�ڱ��>��"����|�.
���m4D��f�76Xb�,��J��� +�MO^�$mۂ~^�,�$]�gs��G;ڱ-
9�3R]?|P�i�N%ciܶ�ģ�H�}bzHC@���u
��	��g��]�.e����y��ݜ��Z5�S0�ҔI�Δ�	 �a�d�����9Ӓĺ�q��uy��,xu�D�� -D]21�C�^G��ƒɱ6��8��~��j�#7$Ώ��#���o�m~%��y�h���n2TqW������Gm��;wlT 6������mN�kK z�rB�|�Cb~+���~!�-�;쒖L��M�o��>}@7+��U#qO[0Ū��&y��Ke3Tsv�5�ke�~8��t�/!�?z5O.D�(�0��!j:���n�h0�5�^�;H�4�]!X*�+q�_LELP����ܫ�:1˥�@ٻs`�Q21����4,�B���b4�'�l�
dX�Ll�����5pYp(�:31��q��ҏK�E�cF��:���NR2�'�?�p�iл�E�m�86E��UX��Z��7���qh��m�'l�cG4xcJ-��;i��}�)��1�k�����Ў�n��n�WF�s ��D�Mr��0�����R�<��Y/l����%.���!z��rۧ�,����"W��L�2TU��e��f9j3K�4��r�C�5�p����}����
����86�X� �}��.vs}�U3�F9�`c�PK��V�W��W�vĪ��s˸ ���Og�c3��:L��ꞇ�;��1i����O���Ƅ���M=IQ��"�O$)B-���hWG����'K����?Z�)�v�ΐq�!��5H�NC6�?fM��G�hDkv�.B�º�.���c�>4��(�#��&[d#FD�a�M����=ŋH#F���C���jbF���Y�� ��8��t�j�_�-��c�z'��$r�蓶ok���c�J!�
�y[�s��#(��?$�&:.�b���//z�S���zv}BY��ޣi`.�9��W/I�qe�[Y*�6�����A�x��ïG��B�܀)*��r�D�uD�wb��װT��ڣ���.)t�.[㓶�h�V�Y�N�ճ������z28T��^�U����^۠H8�*��sB���A>�[���D�a�L6J��Y���5�0��e6�_��Ӣ{)Nqv,��!ݞ�	�E�&y3߁�����R2(t�[�	a�k��K$��-.)��z}8[kX]zǎ�����V^�����ƣ���Vz�:_ K���i�s"�؃��G��Ÿ���8e^K燴Z�A<���ټ#�0�בB}mңh��W�j_����k���[i1ɕ��͵������P�����9�N���&�Ѽ�u�n��|��wѶB]Vn�@	��y��g�Z�?��i���<d6]�|��l��T�Z���loǃ�T_�|��y���W�������_�`����0�qe�^�A%��,EL��<����9�� �b�vNT<*E�/������%1���6ӂM�J"���@��1�S2�����.U/��61�q�E}�'��:��̃��OB�`��[�ZA��]��ɻ��ԇ��
����\� �\%�������G� �@d�.bE��4r*�^6��k��l��+\�� �<�fmV�#��n
p��{P�Ċ:�[b�"��y�)�p�!��Kf��/�C�L�F����%��8�58*ޫ���=Z��Zn����{�K��o9���M�F%*S��-*�R�,VG)^��Dm$eK0_t�pA��+Aj�?|���ؗ8�|ӵ������Ru��2��2䤨�_������@u���D����Si���o�<_��R��rt��Xh�Y�+*�3Q��)[O�s��4o��h�Uz���$�\��*ƸO��K8��7�Tzߖ�TW}~�\�]�Ԟ䧏�ŏ�G/���[���9 ,�����v�ɃX��j'�DLj�n� }���\w��pj�����O֙�Lz#�}[@��aōq�GXl�O�v3A�i�6r<D�i)��4	�\�0�B*��N4n�Rh�a��c^5�+�d9,�2���b��MN@&��L�L�D��W�R^�*��0 �E�Z��@����`�k<���:W�vf1�ϕ�S���h92D�lq��r�Yв)j�L���I�
��Y�[�D	0�-��~ ޢc� ��,j1�9-����5�5yb4_�c�?r�8���~>Z��+ �x�� H~B2k�`j�QZ)���!����#S2�]���M+.��G ��S�n�8F�د�U��
��E�[<��a�1���g���k�qZ�`/���4��n��"ޒ�Ir�{ 4�_~���z=��88�at�VY��r�"��M�懈y�]X�:XZ�Z又��������v�¦��!O
ѝȑq�֧�fWm�[7襅�΀�ƟGmq��4�cl$�\�'�bp����<L�:_;#�߷]]čh�������
���]C��5�f@%[C�MQ^�TEn��L���k4�~H 	��]O@�<H�o�<�v����N"����rޜ �d�f��Oމ�RSVeMLC9����l�A�E�����.D��<x=a}jtud����;�~	��i��]�Թ�6���m�K�����B���zI���aq$܇0̊��}3���%d�a� ��� FK�K�k߅�R;��3eνF����F+
zb�ṞMi$�5�g�#��lt6��Y�e�$	T��5=T���y�6�M>���41u-� N��9%98�7N���Gq>q��,����l;�@�y�'���H�����ZUgs��vٽ��޴[�������	X��}?�s.�8ޢ���bcH�j�F��M𠜧�M=$9U�>n�̥�7/��N�v܍�ىνח��1v�u?���$�5Y���yGȗ,��?m% ��"����g�{����k�!�B���³���+���2����?~�^�|wV���ȼP�JZ���Z1����#Qi�J�%��q��,\��p���2�)�_�Ҕ/V����ùDp_�h���A'�;/"W��6��o���m�r��h�@v�?���d�/ni_���g�%۬��ܳ���C�9���(s�jX�%)�.�K$�W�s�]j�݄\�D�%�= _n��[MB7�xu��O'zi80e�%��2<�Ac�Y�c��.����=�Q�R~]g��ʇW�!���r�VK+ˡ�G�&*�7���R���
 �z������ h��\3�B���FO8*.�	B���!)��wuw�x���ͩ�Cހ�V�7|	M$R5�������=�U� 70(n�Hrm�M��Z���e�!�0FXy���&s믘O�`N ѝ�����7X���0S�1���6�y����fZ^�$YN��C˃ڕ�����	@Lh�E@�DP�τU젠�S�&�'��A�}�7}n�|"�y��z^�1�����#���9�Ga��0:���w�*�a 4ݏ �GE��^���h��t(�.5m'9<�BƗ]��1�uPhq��.�j��Xm4���A���p���M�u,>��41hU��ͯJC̞X�Ͽea���xz{�G(�@��/�������OȱI.u�9'��e@�$^��'�⨳{:%��*��Rބ�I�X�%2Y�U�C��H�01�EnDT�F��=[����������R��mNO��� � �Zvy��C��?>\+��5Ѓ`A��)A���,��Ӏ줻@P�q�]<FA�H��.��"]8��Ҥ"b���$P�|������DrÖty�:�����Ί������S����yn~�u:l�T���o.�6�qQM��#�C��=ٵ.]�VEWz̶���9`�+A�z�>�#�v��h�듇,E(��~cr��9�H�)?����Z�f����id���C���{$y٘�Sr-[��V�*�;�?Q˺��h=w�5Г����hf>~8�j�˳���6����J���=�z2/b�;�����dt>�d�6��?vY���ʕ:
'06yd�и8�ג �՜+y3�������צ�����X���{�b��l��'�iU�-�pZC ���m�ԛboS �7��U�&�!Ȣ��R����:�2������\�7�rV�`�4�%L.)'�aj8[8%Ռo��}>tNW[�X�2��&}�0 ����@C�ʚ���z��[��'8��D�����4�h �L(��R�X�|�����Jd,r��h�2�p�1��Gg� 	�`�#�:&��׵q���Ѱ��K3�}|�3��Z4r{`zˎ=�I/\qC��]p��d��x )G��.�b�)����Ͽ��Sv��i��d[e���S�"�!��~��p�!ek�۩Ck�С�Bˡ_�����:
�H��] רe�����M��8%4v��F��Q!�ޘ��"BW'H ��h�U�ƒ��u��>,N�w���p��՗�Z����֫����Լ�R1�=�0zS�c"pLȫ��U��*����\�.m��>�>f�a�8K"sUA���R(���Q����j:��sA<U�,p�1#�!e˩��ԠD\��h(��dKQG��dL^b�w&cu�;���p~ʸ�J0����j3HO�
�V�'&N!Zȿw��I�Q�G�<��?�oJ!4��'��������§��x�G*,�����;��ț����RZ)�%8Z";���ʱ�eh�A���h��5�~ǘ.ڍ����o+��2U����|�2nG�Ȥ`�	hi��!JFq^|���8p��2@
/_p�<���/�Y ��>��#رSL����e7)}f�ۙ�i�`'У�݁�=v�U�tQ�H���z�������W�̫��h�*t$�<8H���n!�Y'��w��zv<B��o����i����&���ٺ����O9��pvl��]h�z*z�%�c�5sT��}��!P��2遄��+�������!S����^�0��{Hs��3���
3��\�U���G��sd�٭����֨���*$&��|`���ߩzf�f��M/Ī2�B�#yW�O�bqz-x���G���+�~ԒS�Ao��_@��i�ӳl��ٍ�֍Y�_��F�u:�5=��,�Qߧ�Y�a ��N\gAe�UpTp��\��t����o��L-Z?����҄1H�~K�W��k�ύo����{�� >� �N��J�?����<P\��ݐue�>��HS�hѬ�l?�$���RU��9��c@��*��(G�h�me��P���F3a�^�M�|H-%9%�m.5ʴ��Nw}����H)6_���:Ƽ]*�)w����w�L}�X�9�O0���؞(<�,	�������2��I#�kC4c���+��)��>���~k&#����,X{`v>��qUI3K����$2�[��h��l��/Ǩ=`I��d���Va;"�E�fmC�71�f)����*�DE�#�����0A�lw��CF 	t��LOʩ�(�q?�|��F�G�=�Z�:��ӈ�����f��Z� E��w�+
��'����Qo� U��$�(�g�Z�m���=4V��A[��-`;.:�PK�Jcȫs��Om�qiə-�SA?})�X9�q��!i��� �+��~�Z"�H{���4�:9B7z�(������AǉN(����T�"o��
�V���$�tJ�L-��!X]��Tx@���`���5�9hD�S5��;#J�L>IXu�(Sk���;��"6�Zn��e��Yp�
K���l���H�����r���x��"q����Rߦ�s���6�������Eh���`+q���Q�K��k��o����C��]��i�₍z��lgs�%\�n2�P"�����_�na�ƞ(�vM�W�%yH,,S���dY�p���j�e�f�JFs�8r�������?��!�v��t�]���jV�杞�ȸ�D��}�y.��}�zJȷ)eaw�§M��+	�Lt�M�����:/�OM����F�-v�y^�<�n~�:Vw��/Y�ݹ|%�-�`pj�g�׹��v	d	�ӫ��Q^3�ӆqo��B��j}_�"��
�׉���/�r�������ME50RWhߩU�@2Hɔrg	��� ����Xp�on�"Mm߁���=[nk�_U��/{(c�c0\��,�@zt��B��3or��q�
����P?��ڊ�v�� ���u{	�<��������n�Ɵ�ɖy�u��
�)ԁ%Jߊ�^�9�zCG:6&bUh
��p�O����5F��҈��Ar_�-��%p�P��]�gu�䞶�Ԧ��*CF���ס���$�btM`���;'l�B����B{O+��2Q�ap�̋7:&�t6����$
��n����r�jC�R}�E��7NǑ��aTyk�*��������H%a!���H �-l�2��K�����m��3~�R�	�nZd��b��J�M9ZF��.�
#L�0�c�h/���މ@*�zTm.ൠ��v��"XWU�:,�o��w�F�+�M<��w�����
/���SƯ���"Ԍ��8�>����8^x��z7<!�� �W��>v%�jm�f�	�W5�қ��QH�:���5�%�`A�=��}��W�#F�
;�S�\S�]�@u����\F/���4PGB�tC{�*����?N�S�󕻺�B�'NՋ�1$���C	�n���8�JO��׀q>얨N%2#YJ^�,1��S,��K�y+H����T<�	�c��N\�bU�7��f���ݔ��@b�eN�S��K�3|&1=w����륳�ML�*3�|&��@J�m�����&8�x~Z����IQ�\v�#G:e\:�%�`���Tl0c��(�U���Da��1��HȠ�dR�k@M�Oh�ڢd�mh@j�$J\����.V���L�K�r�Jtu�z�j������Q_��BWICO!���`_�4�h^k���%+W0c��f��t�1\1��n�ٖ?�4�Ey���]�n��:�0��}: �ZCVޛ��3=�ڷr��`li�$�]�*Ҹ���"�{H}ωjw����]?�4������0��M���N�_ץ�k��k^����� Ȉ�K�������|5�_��[��|+�}2����〇�\|Ő�f���ݮ�5l�3�1�4�/�����9f�c�C�������'��?�����B1���rr�> ݵ-���',��^���D�\,D+KO�878�� `����3/�k��~��撃�/25z�f�,���H94�����a�����p�8L`�|-�8e%�������O�f�Y�Q�#�'��Ifv�$��9��گ�(�=M��'�G}%�۳����h$�# ��*+��Z��s�bU9Լ��������w0@��0&>Kn}�\�ٞ����B:%���9���3>���@� nt�� ��U忈q���|� ���_���j:E1f����6ػ�	����O�0��.t�U���C����пAzF�lE4AK�$�=<*{�PQ��l�nr�[e��5M$W��>��؇�
ưa0D����{�[FN�z6Ya�X�`a�m6#CL�dI䅖���2��k?0EJ�(���)߭�9=��T�+`�'��_H�!٘~t��+
Z�xXk�?��X� �U`Mz�Y����4�*�����ֽ4*���&�1QZ�J&�
��i�_\���X�rL���ޘ��mT>��S6�:�?+�����YD�/��ȿ�6�K�K�Jfɤq��������Mz�GE?�dz�1�M�Fl�_�D%�����g1Ֆa)�������j�_R|�{�nW���I������r�.p��X�ah��|���
]�P@_�4��S�R�����{�M&�tBo�y}��M���ŷ��?e�*쑠�z/�t,�a��R����d\�ť���X~ۉ0���a~���qՂ�{$��X��kL��u�*�����Y]��G����4����w�f��z|
:mK>�S�ΰ��� ����&�k�2�5JѼ�´ׂ41x#
Q�xw���i�W���N� ���q���pL��#�_4�O�͡�6)�F�Yf=D)��Z*lZ��@J��_.Ǧ�B���@�7�\g�dm\�����%Vh�)�/қY�Z �.�^&���j.0�KsLK[�"��w�JM!ӹ���d	�T�]���n��P��E����N���u?�p�q�ҾB���д��©�&iN��]��h��i�1O&�0�}�v2��s1�$�g��
`ӥM��
�o)/�7Z��BSG*�L�Œ�dE��v�]٣[bE���$I��Z��a��_�|=�Eҧ�v����{�{����kC߮g�f����]��pؘ�Ւ��2�R<����(l��{G�NWm�̹AD #���Y�����FT�z@���H�l�r���Dm�3A�����ֈ*��Mo�Uu�� �֚{u���(���p�X&�~� ���k�-4Ս����h��R��b}��:1�#�R�1�@�W�e��}	aY*��%��魥�U�5t�d�V=-馬G{�S�C�̰�Ћ�a�k{�r��^��u��?#�Jv�,_K̹���x�avn �~��t�CȞ��>���6���'�%�2l[0��hWP�@R���ķXO�s<��7��.>�v�dP����!�ŋ5 ŕ�Qtn0D��J�xY]^	�<�_^�Rc^�m�!!l�S&��o��C�.u�܍A��$Z��%��f����1eѫ��e=N�@���*�J��H��\�؏J��)7Y[:1
]|���Rq�G�8
�sߺ�@��x	;�]k�kd�k0cS�L�?�$��0E�8F��гGl K'v��3�㿊���GJr!=L��w._��qICwO5�0��O*�<e�Y�r��ķ|�[a�Z�s����8�C;�e����S��-�nQY�m��%�+yV�����5�)�_��oW���r���n��f�I��*�ϐ�X���|�c!bK��J��4���!TXn��=з�6��H��fy2ў]!u��5��Gx�5�1� ����$�?]�{z]�+��]HF$�3X	�"&_��%�\S�!�A8[aۯy����^�Ru��{��ĠP��|���5�bRJ�:�=�,A]��l�N�ٷ�1��v��n5O�f�\01YyE_�@-�ֿ?uJ���g���mɾ(	%�,�l����-�ipG���G�cM�ʇb�DCd}l>}ʠ�z���U!��Zv)�<Fq=�]Z�R�P��Y�</�]J˼�$�����̊Xv
�O�Ż^�A}���#�D�X]�5���<�"䌵nԏS�ߪ>��|��5�JBc[.�VTxRu
j~>���)���
��{O+�~@�G���R(x��za�Ȓ�I��s7>��m$@�%CN|m��;|7��5��pG����v	���3�"�[Vo;Гl�^��C1�9e8}3{�S[?zX���Q&���a��%,߈�r���]ڙ�D�@�M�W=R`�0���ɩ�Û�,A-�/ r��nMd��;��U�W�Cf`�{�3V�M���~�U9�`�=��h'elwy2a��{�ᅓ���0����kjs���+�-ǎmZ;�_�%(]���˿g��ó�s' ��b �2z �q�ҙw�*�;>��ڬ@6����\�l��>:��ԁk:h&�&J��hb���p\b����F-�#-�2>�^����p�+h
�����C���nrH�yB"��g �vw��T���'��6�����e:�8WRD�C�D���N����pk�����?�5��T��D��ٰ�?ݩ����E+
�Z_(�����8�����=�+M̈́�X x�?IT�MSF�s�EZ�4B$�s��'���Y����t��Ő�
�����YI�DV2<���.�6ޒ}a~C�u+��Į)�����C�Qc�. ��0��3qS��D���;~�l�-_]�i��Tk�)ò4(�ܕ�s�Y����L���>����p�9���v_'z1�}ȜC�M�er�iQ�sۗA^��w ����I����/�����Gʖ6�]tF�(�RKN��6����2�Yx^�I� *�V����{�|ϥ	,�N,�Z��3=��7
�s�&�]� 6�QM�=)�V�6��-��s�U���Ǖw,k�Kܽ%w1�}�O1�ѿå����J�5�h�,u�O���*.i3����r.ʰ7�އ�2��!���b��ZY�CU�q�8HᅅFCR���TT+���p��͑�ܶ�jLS�6`�`�l�%���գ�;��1����e@Ȳ��韢�������=Ui�0����f��5T;����b��Z�ߖ���oì��a��f�z��.�r�M�Z�*�Y�yI~) �ԑ��'^)״� '[��=qMq0Cm�!��YŃ50�~p v���i}.4&���Q��6*q�͋� �����FV���V����>���oQ�/�C,a�Ҭ�� �#�<�x��Y�|��{l�%n�n
аS�wۘ�xx(�.j�'���Ԅ�!�EH<'��aI����+, ����r٘��"!}(�~	ß���S
�9,$o�GD�4����y琱��>�7����Įy,#I�$�����/�_�F���
4�7Ha��3`�؈�?�I�NE�:l�k[��ā��ݝ��n����~��f�"��t�'�|��D�t��@>�y��y�ǽ/;�wC��B�.h�~�\t˅+�4�`(��������f�Ă����;�"�.Nvz��o�2����/�/�9��ѷw��ˁ���[&�{/���M~sKr�����3���i�-�d�}5�F�]Ǟ(����oN���1)����M��ނ(�@��%��I�i-�����k��2��I�"�uT��w8�:g�32=��Oͪ���?Imؠ��M g�����k,WIs�L%O6� ��r�?Ԍo噸'��^ T'{,�*N(樣��S��a��|���)���bJ��7DÀr���ak=�Aߑ�y�.�������`oK��7�@�e)g.��f��}0B�Hf�?������� �5l�-�X#�Y�{/9+/�o�}/1u��#3Պ�95���Ӑ�?C�h�9��r֭턈��i���;S�-i�l���y^m")��kO��(z',�k�E�k�z���j��z�3#U)�O��Q�A0jc�
��X�����qlNV�"�±H�窱��SE�k�ˁDlj�:�4��α�&�l�2)���*�=��r�'D`�[�
��а[o�2>ئ�c�H��HǓ�P��RD�PC�g����qZ�QW^��[[Ke������@ӿ.�ʀ��ʕ��K��@0i��Z"�S�ڐ<.[�Jk���&DJ���7`u`��%�<��X�\!��TL	H�"�.?�����������<=t�Xk�􋉭��H��ʌ��mȊ,y���x�D�9t�t�r����c3���YԸMY�v��9c�lfr�@���Y�)G_��@}R5�Z�%����G���'}���SIj^{�lO��V�d�ޙ$�|��
f������"��=�B*b��N?�o��fũP_�!�T��&�	�P���wu�q�6̵y��Y�+NFW�{5MU��?r�ˈ����t�*)ERk�����E�����@q�&�rФu��
�� S +9͚�����!��ű^�:��"�Q\��^ �z�"�Рسs�^S�@B��z���;�<��6H���MS��|�����:v-��s���t&?J	k��|�A��_�.��=�����������La'���b�ߜ��V��/y�kI��A0�#��#�3W��%��*Z֥}�U�=�No��_�rj��2�L�v��\��3���7#F���:Q�/ѩ���6���~� kB��0�(Ƙy"n������IcU�!�k>5$�he ��h�[&�� T*M��4BE�u��׹�4o�^�K0H:�ڪ��BC�p�U|�cP�/��F���`BJR���g��ʑ�K���#��ZC���l#b*�r1��;�Kl�g��1��s��m�������L�l)8ÂF͜f	��"EG(˨�3���F�Yr��&�7FH���n��见�����C�+��I2o���U��q�g�����%�ۤ�>��p�Ń9�����歍ړ�?4��L���7h�,ډ���!�'�}*H4��l�����/�{�S4Po�o�e<�@7�+1:_��bg�:d�*��Pne��K� S���n�0c1�-A����W��3&�`�<��yU�Y"�-_
��O�G]�lk�ħK���A����5�5F�yt.���G���c�ס�!yN����"ު�>��I��k,�/z{e�?,b��#�n{�����nr��zoZ� ���]���	g��D?j�y�������	�<q��Ժv�|Q�Du��F|�|��v�����5]����� ͐v�=�!����,B��^S5�4��~�����@�_��5|�v�A�0r``7�]C�"8t"���dE$�����.sh�:+�qͻ��3�E��8"
l&��	�JB�ʋ;3��@�@�'~ɟ���P��]37mn��G����0�%ͬ���>v/S�)��6i�V~5�bP���N���J����z�Ա#{������k#Α��LYa�P4��=2%���"�tX�e��I����6{�^��x%9���̴���F�)�t�P�WJ籾��(�ϳ̰8�%;�����qN�4�cDv�|���(4UG��:�u
�sJ�R\�Tݹ!'�`�Y��Ҧ�S��_O����5�f>��I�+��C(�7,���G滾2���a2����X)8��"y��*��d���s����k�"&׋��ǋ�4���VԋC�hK����x!��վ� 5���"�ݴ�@�SkL;�^���2q���s'\���H"�͇�����RI�@]F�����}�P.*4���{;'ꙟ2*M���3K��:��p�*��|��8�%iұ�V �.�%.��rc��� ���V��7i����ivQzKL�)�;���<ٸ��:��q6}6��i�k���8�ϣ5S4a��k�(���D,K"YaSD�'�
7�/�UL�_��n:���	0�l����t�T�zY��3��ۮ�E�����m�S/H\]�f�o�g�ua�@���XHw��[{������LK�u�}.T���6� L�O1GR
��^�꫇�r6���c0lYQgcH��c�5��}g	���zZ�'�vL �&�;�w���F�6"�Z�ǚߛ��#��6�J\ڤ��,Nk�e�r"K���+($�����>j
���� �S�h[�9�;���/ơ� ����{�.�+�h�ӵ#GYS����ˣ�������[3��V5n��S7~)0�Z������i�M}�h):�	^A��Z���kZ:i�zSAR�NK��zA>�тn�&�����ֵ���xܣ�ұ,ng�f�J'���["��'���"O�}B�l�bhX�(�]����'��3�)�gQ%��<f�K�fI��X��?ϕ2j��P����b��[vӛ���{3��9���MD���6���G��p���ܲ��X�W��_�o�.�i(�2�t�#���dH�.꼲��,��� �O�L�۴�#@p�X^ctJ,�?����Gg�Bq������R=Q$H4�q�R�oƹ�Ÿfz�c�g߃�s��پ ���I�-s��c���9�ϥ%S�$7VK(Ů��ng��#0s}@�:�i���P ��8�H��K�4���v*�q܍1T��6@(Q߸��p���xu�J��'�6l���pg�^y�B������������D�/�֎�=/ҚLզ�,�Y�#�G��8f>N���ӡb��Iv�Q�8��_کd�E=!��D5&!ߵ�L�1���9��X|��H���]Q� Mڂ��$H�_	ż� ����2��v��;�ߝ>Z����ƿ�0eϮ>��\U#:$h�ă���}���;ww��?�@*�y�iI��,���j��'�W���_��}����q�_�"~�z�G&�#����.�ߌ�H�Bn�6no�H�T���[
�]4j�u:}r�k̾o�����T�^i�~��!a"��!��i%I+���"ɧ~�R��PnÅ���~ �^W��MZ�{��P��!9���PU�}9�59�?E�_N�(�~�5��{��aB���:�#LS;Ћe�6�f�l������)p�P��"2�c7�`�wM�{�!�!f&��y�{�$�0�L "���k��������}�r�*��i��f�EFK��#lڄ��I���j=��s ��}�sc�Q��|�^oz�Ql����"��6D��s��ME<+�d��*L�/w{w7ۆX�op��݊�R��]�ph�P�eap�z���G���t���=}��n��wM���j�����dn��Z����b�o��],$����E���^�I�` ��(��:y�h��A�5֠Ij�E}��K�����Ge}C��8�8��(��n"���DyQmu���˷���M�c����ܘJR�l�������R�'U����d�	�6�A��r�p�Z-�̋/�[����r"�Ǖ#���h��n�����z+���gWϫ�a�L1������a!sԖ}���oH�Ӆ���i�]�3���ZMs�a�)x���(^��z���@n�h�
P�G4�<���t~�j����|I�I$[�\؅C�`HPaN�1��ު�6�]�~U���o:�� ���ځ�p��v+�M�q�����YM��м����Û�v�4��y��4)�q/�M���K��(��~�{E�H�Vх�3Em���9�^z����J�y�2�؏���'�I&�L�ٮ0(�=�ӣ���L͔��`	��D�{ dŅ�Z�1/wF:�F�)�v���o���V&xJ�)'�Nfe8���QВ4Õ��k2ܞ=�wm-��>> �-��H�av�2_��*7M~3s�A�3��9���$_]��P���m8��87q���豅M�����?�à�C�AGC��?^�kam���w� �+��e�
��H�P���j����*>��}1��,�X"����o��z��0T:�'�3���/6F�o�\��aPz˖K��M%A	^�(�=F_����0�'�I3��T���Hmd����Ȋ��u���3��4Ʋ�^�1���Gj������xS=�����`�4NC���� zZ��V�f�?��~��ދpt��ƕeu�:�#�7O�mO�2a^さR b�jm.��Qp���2Qu��L/�q�߁M2��g�W�!������=zQg�g��Nb�.�L�/!n=��]�;��"��}���<}*i�`%xƤCW�SrV�g�>s-z,%���[Rx sT[���ҿ[h��);��z�Q�=ip=�n��w���>��؍R
��#�W�uH����GLwLN��D ������(Ru�8,�ʌ��8IcP��4!�i�2�ыNk��m�B��d".��Re�6�+�3/�X��4���sQa��b9&شtc6m�6��όkDU��W�_���>]�����L;�i]��g�XI-��L�ܮM`_���\)�{�}%;D��Z�״GT1�yΙ����"��7o�{�h��k�&��.��6)I*}�-#{.q��R�ϙaSr7?�s,��9�|N�I��:��7*9$����>Pz o?���=&����7�9���_&�����+�+�R��hs�J�`�8$�Gp4`R�!����$�9��ˑ6M�/|Y9��C֝Z���le@�m�����-�1w��91%���l�-S���+X>��f�_G�'�ԌYxą�ZF�)�L6��փz/�"MLB�$�K�����B����8�|�ǯ��‱��x7��>�P{�G�*Ri��3�#���ֻ�K!�?/tM�E���ˈN �'�:��T��ҝSa�-��-�3	� pb�k<̫ܨ�7;�+�ZG|�	�)8�C-��B���i!�#bb$_,��3F̥�3'���;�FD�1/�toc��ܸZF�Y���R� 0�s����;$I(l_�x7�BlZ�V�!���"8��F�Ŷ���mk���*�bg��ׇ�,!���	�	�3H�5Ë�}u�#K�#���>���nY��V���ߊJc9�h���A%�T$�Q�-�0���Wv��Z���ߒ㋹�?u��g��Q�iB����Z!���a�P�%�K-�GVd9��ě^�W1y�1��ş!~�Zx�eԷ_j�k
��4�jy'�q/./�w���0t#Q�{�@7NJ{���*��d�q+2l���0;Zb�޺���B32���� �}��}�f��i1N���Ë�%��ܽ��<m=�D����u����_Du���X���(��,��#tG��٦��~^���/�J��a�����1�{�"�ZWyjW���b�
�u�>��X��0�&?���T�D���l2�?��g��¼Xi$�lZh�f�f)8�v+��#N^��Óm�{X�M|?���kM��=��Y���M�#����^ct5���^��!Ƈ�(�9����g�j�c's�7��"(�*�TM[�mN���%���7G����[����� ����y�,wN1���`�(�K�]��Z	�(#��N��Ç�c���Ț����}����wP�Ǡڥ3��2��� W+��щ�*mCg��f�ҋ��Y��3���Ea@N�,@�1��*���
�+�4����ݟb�]�+����,����)�l��U.��Z�l"A�C�޵��佂�Y�7���l��W�����oyn+5�F��H} ��oS�˾,�Iy���51�hĢ;����BG���Q�K%*�^Z�\k�����F�g��v�f~}�=��q��i]�����)�V5��?Ԝ�T#�=�"Fb��J�M���k��`������$�5��GR�x"��������.[d:#E���K��]"� +�#;Wr�R�NR$2�p�c�[h������ʲ��ߺ���ث�J=p���i�;g} �<��:�<�g��?9H��^d����'������p9*�fP!6�b��˄)������[��!��S ����6�$@��S>?���C�s�(qC_�E�6-v6��˚�ڇ�:M�eh�>Y�[| ��bl���<23��85!�'���r����<R'�XE���ٷ��a�}|��n`��a��s�MiH�tSdc;�IÜ<�ȅ���RM>���j�?�=?7�?�Ĵ�d>�<w ���~�D��Rl�	��.�I��n�+ߘI��z'w��}��F�=��M���*K�1�|G��	�'��/oFhU��������8�dç?�z���Ux�rT�lZJ�Gq��qML��1/+��N��Z�kv��,V!��#ST��"���	��t�~�Du��p����ʚ�?�{sǣ�չ'z�v� �5z����T��'��yЌv|�[@�V�E�j3=3�U�������'̝�s���iU������B=���pu���!������/�q���*Fn� ��FNc밗T�dA�9*�D��_�!jH|'n��i��["���q������-�4��Z��Wϱ���V�Ǚ�-��✹�BhdQ�=����p@"�B�֛��.ˑ_�ș�1I6WV�����-�<tp�R�S�y���D��O�������KM�^��#�]�Ƶ,�O��i�ԡC�Q,d�c��^��*�B��f�zZo#�Pu����5��N���1�������ϲ̓���'xs�7͍���fN���3Y��#���W`�xd�
�6��	��?�>v�=
���v�xD��;ˇ��uN.�!B�1�b68�>L�Jd�}��?�4�G�̶��!D�ԊwZb��L�K�X�=	ߞ�|��&|�~1)�ڽ�!f�h����;1�]իz����@ B�������+�����Ǒ�4_p��u7"�惘��[�R��D�	Z�_�q�Da�w���)��u�!5��0qo��AG��Gӂ��`/�-�[u��.�,��þ�Qy����(�Q ���:�5���f�N����ϳ#;�M�Hb���Jl8T9�[��MZu`41� �>v���W�V�ⷻJ�NǪOfyI{�@�[��o5t�}���L�k��'W�Յ�B�������1����wرq�U�v��,�i��r��,�x��,YU56=!��
T��I�$��iB�J�x���C�.z��g����ߌ��ZL`5ԞrnQ rl~�}-.��A�����d���]8�'���҈H��I��7�V�㥴�1�ǒq�L:SRe�*`�^7I�j��� ��*�E)2L�=���/?*hJ�9[�w�9v��G|14>P=�� �\�#�gՠ_��g�ݘ����'"G{B������	�7�t���� TC7�Q"˞�Leó�7��7�y���b������~.�҉8�%�C*	�4Āܿ�	J�f����Bzq�!X#8XG"{�u����L�m?���=[�dr�t�4{N�T�2�*���ߎR�@��⡃�朇����:�;�$t�S��2cX�0�4Q���(ޛ��ǄG�-����x�~,�8�a��pQ���"����~����8�G>sk���x[��2��/%����Z�N�(��2!���j���'T�ӊ3�UfV��^|��������7.�N��}��B�,���<��#'���M�ϝW�ӬƤ6JVF�\Z���X������z  �x��~ې$��,� �֛f2�;����O'�q{~^�����5j�0-hp��M�z�����} �ݺI9g,��.���f�E0�G��-+mk-�T
&e��Qe����4�v����{�[>��>���W�1�eD� ��F��VǢHk�=P�_��}=dL�Z��eW��B��ٳiK{�'�c&�����iz#�a��u�S*8���\c�ྸ�m �U��dZ�?��4����x%�lȚ 0J����|��+y����ȩA�H_.l�M�c��uT�|�I�k4�
c>�Ț+يR�ޭ��Z@R"���ק'��w�,VHE������	��e��Ћ:�Lk��H��Gn��q�4NK�ʘ�ЍV�V��������'�D�ɮ|�$�����z�c�_^�<w2J��<Oz�9�g��G�p��
��J�isR�8�ᐏP+J?��>��^霷���f���aT�������r^�$��ǏS���)�M4Co����`��
��ү_�I8��Z���7j�?0T["C���	�����c����I�����mU�n:�O�ʏ�-4Aa��.ˉ�V�܋`�[XQ&Z��@����"Q8jk��#-=(�{�&Ypf�BP泱J�j�4	�\�U������K9CL�����Y��A;擮;�N�e�",u͎�Qb̺8Ќ��{�� ����7�mȪ�ځ�� T���7�ԇ9ab3�2�C]@� ���7�� ;	�_
"Zq�����Y�!m8� �{\[�Ͱ�4��B�|� i��LF����I򔡿�3%�d��t��k�D���=��� �ޒ0�낝@�c)Q�,�m�����(��B�z:�n�Y�Xq.8�<r%�n�ǹ.{!b�6����t�(U���!��	baLv4�"6��,�D��=L\.�����B�26�e(>}��&M�g޳A�i�z�㦕�K;�Y���3((�9$��rqN�S���Q#����&��;�^O\�����n�j�&y����IB��lj{͔��wVQ�E<� 9�rw^��'m��@E��m�YY��S' ��?KS�b��`��x�O�nK{0�yOyo����;�E#.]A-�t� �e�=�3�F殈g�e��ߚ0�:p��(X�f�9ȧ�BSz����:xv�1�̶x�<}�s�yd1�'F�O2����D��_j�:�!�AJ�L�n	n���O�G#���җaz�Q@�xu�]/^R�]��p�d�A��a�jk����6[Num�К��xڟ���e�k��p5��|�6r�D�K�6 і�"��1ք�3��-��K�i���[��D��ޟe���'�2����nJQ�Yk
 �28
��2a)5���>�9�{�=��#"�_��p��Q��ꪸ���r狑�.`��Am��a��[�JJY�5�g<��,���)q��j�E@�-���D�Ѭ�	X<��j�RH���	�W�6�Uf
��nN��ͩ<p
h}�v�R���r�ƽ��̖�����8K\�ԉ���=����0en�r����3����>gg=��6�~|���l�����L-�5���N�,B��� Iq�8�b�Qg��l�8�qA�����i��_o\�@ޗvm�}{�MCF��i)�`L;�/Of�"?��TM��1��q�s=絫�r�%�Y�~J8E*���������g��lP��w&r��|�)���"�|*w�Cz _��AH״]b@�C;d���$�z�1�Q�383�ǰiE9���7i��z.�'5�����$T;Cd��,VB���j:x:��<�pW�n@BlS�����\ì�X`7~�.wc���J"ߖ:?6�O�:L�'�;���H��LY�ن��/�~~M� J��k�?�\*�Wa��Qi���0� >����� U��"S>�>D��(CAE1�}�a�&)��-�0ߛ�G+�L����F�޻6����w�\M����"GC4c��A���Ƶ�q�Lpn9
v���T��I�0�H62x��e�@�K�D_�]+�(�]<P\4��Ь��r�,o�uP����$�| ��<�I/�c0J��*�K|]nc8^)A�)�n��$��{^B��Q>�*P���U�W��Qr��iǸ���O�k�7�H���1Fe��9.�V���gdF�HZ��:'D{���8u���eV��=v���`0�Ϳ�R0�j�iA����Ǩ����(3�bO�'E������2���b�@�vY��G��,gGf��h��W�����L��Be�0� qo��֞I2 �R�qATi-SrO�ua�IM$"�מ'%�"�!F�����H�p�V�?6����`���^'�Ő�7V�'�y:���j	�0~����	���S)��Ў��&U�kqh'���@��"uCn�[�*K�� �V�7�V}黨���o�aX��0c:�A�������^}l\�xɰq^�v��B�%R*е=�ք�T�7�®D�~�N��ߊϜ�;����(��f/�"���4x�s������0(��k&������P@䀴��&��nR�2�L��+���J2��;(μC0�ԣp叿���;l�@�ό+Y)ۇ�9�7��Bpj�K�-
҃�,0�ו�>�od�w8%�Q�s<3���{��_Խ�>�evf�w��Ҝе�:Bo�P4�B��h��U���<���8��/���F��c��S-�v0_,t#�L�NkK�$�H~?	����6�7�E��
�և�a���s-�;���|�T ��"*
�`���vo�`9����ɶP�ˡ�j(����M ���!"�ί�-o.�4/oE�3�FL�"��K�1�/{l�G]	;Q��0CQF>�Y�q�@��T��N2��	'7��'?��8ʗZl�(��BfW,�K�n��G͛��:3h�{�� ��hD���9�?iEĶAؚu#;�-����儱
D�?.����g�)��iĝf(�"<\�j���[���MV�u�C�]pװ�[��0�Q	(�مu��x�q��J�f��O~{ji�+�����{SޓEMx�_�K�}���w���D���0��j�
�gZ��n�`%� �M�nȍF�;�$��n[��-0��$��9Q<�)����F����F����Ҷ/Vj�S?q.ǭ&ׅ�����m�ĬH烿|����d���(�;�����Ҵ��#@������W���D�Ԡ��
�����4�۽#�:��KA�'����=2��o�����&~���3�RI��F1s `�G��мG� ��M��"]a�*�U1?�����\�M%���N4��,�5�>�c�)ldc�৒n����fBT�i�g}Cs��h�C,�P2��;QS`
����f�9��J�Tg��a��7�>QU�x�0:G���i�%��g-��Yj��`�b-��Hl@-}w���L"�$Tވ� �!23�Gs2yFYr I��9Z"i����5R9�4��"��)P�씵3�5C��N\��Z�?Ȭ[���}�<�! S����c� \08ijˤaL�V�Ma���0bQ���{����sκ�~ȧ��#���W�[u%�5GF�.��.������ML%��E��g�e/d��˦��T���]�����n��pEr
ɸ�g���W7�YyT�!�*�̅��9?B��,����i���5y	�>n�e��o�����A�J)AI�U���(�HPe��<����?�ƚ��B���������Z��g�>[?p� \��$�H�>Co&�㜆%M�=еp�VZ��\q��ď>K8�;ڸ�W���w�)��o� |��D��FV�4Q���{UR]�9���a�TU�5 \:u!����hϙ��(���A�5X��A]����-^w6i-;�z�. tr��n�g�az�j�*��5M�Y��#����<���^gV���Y����b��8ך\���Ks����Ɗ����dy�qҊ�0�{���M�#� ���#�;|Z���Gun��� �����^ɛ3�T���K��f0*�G�b8�&�j��T���Sz���;�/�fJ�A�l�X��+�J��c��^�
�Vt��D�з10#hH*��Q�]
oa~ɸ�����0�c�E�`�ZÃ1l�����K�2�>�ߓ��so�ǂ�V�R��T�5��8qtJ%������=�MO+���y��7�D
�M�5=_yxH�ٽf�v���ܬ͍P;�]&[�v�jE�C��m��tWx�[��1A]�Y����(�hY��]�p�&Kjt/��r��f�6��[J��=�ԞQfw�BT�)֧�w�[<-`��:�`�H�mK�֣���^5AF�zJ�n6��m�����j(��">f��Y�����sRj�B�e�D��dt�3 ���kaC��A&/�К�pJ���&tN�L�E�n�A9}��z��ߓ�7,+�e����
���  �@PR�᱔�����q�b�l��]���AΞ����4��)���J�t5�u�@���Hf�h��\�{�������解�BB^]qO�����^�X���{3�B!	�r爱��V�Dl���X �P�;��H?" �7� �!M�M"���ߑ�W�u?@���PQ�l����5������~*�Wn��X P�8�dr�vB�e�5��#�����~�L)]����$:Y{w�gj��}�H\l����G;����$u�3�=�����]�P4�G`���'���W����?_�J��4�WRn�u5+�jGA�n�mT�y�ò��]ן���~3���e�_��R1u4�{C%e��oM(��A�[ud�V��.�����+�u+���2a�|5Y�|��컰_��53�u�{	��Rk{��]IS�l�d�i��{�vӠ��w��ӽT|9����#V�SE�~�8�ʺ�X畯��q�=͸��a�;so��e�*|�KCh�Z|��Q�j�4� ��,�Ə8��<�s޺ ӛ�g�`Z~f�$r����4<6;������X �Ut�}�=���������&LA�<�M�i�ܩ۵E�f�j��ty�J�!~:5 �%���W�黱�;�hU{:U~6���is"�zNhZ@�/�)H������cѕ-���,n�gN���#� �����I��^�z���<��0bs��?0Õxh�S�|�f��G�2�>���{#g�/�_�ɖF2���(�Ϸ;!7�I�De}�Ԕ�Զ�`��01a�\��AR�A̞���a7�g��,��埥(���"̇ �u�rB�Kp��|��H�V��.t�AY��m�`<��Q����B�a���»�-[T��m+��`NHEz�J_��i�Dx�+E"l�cYB�E���*�?�N��2�2�\�[�k�%֝ �ʵf�1"'_�7��Z�� �7 ��=�Dp�m�h����;cw���sA[f��pLj~n���t�ID��MV�Ue�r�l��*
pkn�s����y�ï�ݦa�n�~�H��۶˒�r��魾l���_�DP绸�_���4�"?5l�k[�l���:�!`�-k�F�1�nM|0��n��Ԋq�"OL/�:�=�خ�vEj�";ߍ�T�@"O�� �[@H�!�(���&*܊G��++ص-2D�T���J_H+G��{z<�ܔ�qܓ��\]��ifB��(�Vy�q8�+:ñ?LO��E*��䦫՜��𜄪B��l����Б��n4���O_���$��%A;B^��I���oa,���(���+���1Pf�?GY_�iy���k�X�]f��?��uk9��rߟmN@ 'w���/���� U����N�h׋�.P���θփYJ��񥍛AC�7�.����#>u����]�y.g�6O���I��'�{A7��*�C�7r�{d�C�� ��X4�ER�pe^�9�ߌX�S(���Y�Ղ���=�֋|B�|jw�4r��������5�����`�.R-�bl�� ��1�]������t<�����qv�����[�� ��t��b���ì�-�Oo|�Y{$�cNR)i$V���μ��[�&�Mi/��^��)�����?ҔYb+���FףK08�d�n��`���)���1q�8��.�I�Q�5�n��_6)�M�#�k�=���2�/��{�@���� ���9���i�E�� �-�C槹�'��lP 5��b�i!�Ț��ܳs[�]=�zε��}���v�����ǯ(\:<���������6�����3r�n��k�F��/���3 !y�Ӏː�24���`�ڳ�U�8�<� �U�0�5{:�8-'�YT �A-)�G���A�J�|��|�v<Is�c�z�t��RJn�j��U㭦�ᅸI{C�}��(��s�6w�H��O�^DDB�I�6-���>�≏�m[0��ۈ�	���x�b���_���,˔����T��L��d}U!ۢ��<�六#�Ϸ�	�,w�F`e�)�*��'�+���k�:���-fT�Ƨ�P�ڷ��%�&bed�������~}��"&�/����g[8�C�U�U$jk:I�q�|�k D?S1�v��c�C���pa�Q_�3t����O�4��3'��Q�D��;� ڱZ�++ut�D>0�N�>��[�;�D(2�Gu�ZK��'oE�.,��?���V���m������e9G�;��d*��|�%-A�[#�ǝ���-������q�<.�3�DJ�l=�b[�q»�Ӗ��$U��
j'}6��]����,=���)�
�+z�m�2c�-�J��P�� 7�e�9W�PF
T{��`��0贋�O�t{g�l���ȹ���j�6��>� ˎn�����E����v=�S'32�n��{c�� �`�<���s+�)l�*?�0�=4̶0~�	z8P����6&J���+'����Vc�)Yr�w30.I�a*�nV�A�[������¡r*�{Ժ���AoC��� %�B�L�l?�}�d�Tȱ��8�_LP�9O�gm/�5�[Ԭ�U=�l+��b�)��tF�(	����`|Z��X;�cȾc�c�S�_�]W�s��G�%����{�M�-ay��Q�� <��7׻^�Z�����(��	&���s)p��z�r���\��T�j)��dŝF)]O��F�J׶�!7�G0�y({�e�8_h�����<*��ROa��X{���_(D+�߲nO���``�?SR]���[�!�y����;A߷��q�i�v�����U](�����!�t4Z����d�8�0Н9칕7/G̦M��,q����շPS�ogE���?�R�ܓ��_�\�c���s�ˊ��#>`��L�G�m2eՉ�"���Ԍ`7,�:�rǏ
[cT�������s:U�E�G\�5%ؕ�YĪ׺Z50�l	��V�� ��+�I�=�m���O�?q��:ٶ����W6z�AW����9m�D
݌�:m.��;,�gS�[AJc�+��X��76\�{�xS+=UB�����brS72Fo�9<��"$�	�|0����N�(*���<�nQ[�-��x��-]�������cP��<�&�y����Q^��=�1�K|�b�Y�L��fxO&���qg��%�9cδߑ��Bo��?������Ze�W�Х��G&��`����i�k�.̮a�݉43[s�J9AW�
��&�U�W�\[�Wu��q�h�o���5���kp�`P�}�ܞ��U���`�0�� �O�&M�Th���ދޡ�|�����:\w9�K��$8�j+�� Q��7rIn89�����?������#Pl��}o+���/�z���~�Hk\��	� ��G���saOˊ�>1�$~p	����Rں�Jw�fh�RDgq"���;~������D�[�+����2�;��c�M(�G�A7+	%�Z<�/�~	lz�;R��с����{�Q��;�ߒM->bL�Dw�x��sby��e���Y������7�X0kd���3��޷H�ǧf� �1��ü��\UFi��!�	���RR i����C�xt�e�THR:�6�lz��.OĆ���x��oטGx���KF�Ӈ��鶠Ձ貯��H<-�#
6��#� ��BgHaFD��!:�|#�k�����/����|���D��{K��G˛� WT��Z*�4������Nx�M��7��pQz�I���\���q� O�̸[2 �C�W�;����f&�Bs�>���	���`X�*$̉s!�N0�����̧�ٺ��B_��w�	�g��yr[��*%���X���?[�ΪT R�*(MǇj� :���\A�ېr��B>H��2�}��@� 4)�^��;!;u�6�g�oЕ���/<ߦ� z�0ɗm��bk���(Hs��o�r���ϖe��}�L�/a���jl��3���(��L��F!��/��b�Yk��A>��hj��ԃƃR����n�r*�Ed������jN[��@��.��"�4%��&�K����ύ3�B��vh�D�>�FOM��44[��e�/#�85�>����v^W�]̬��XQ)��3�\J���a�a'{5�q�6���{V���)���a���2��� v�u�O��O��n�����#@�su�6��`|�}ΰzՎb���R$#�f�B��f���IO+��@�m_k@5��v��6���D���|�5�UN]����"�X$�8$���b�*u�)M�cO�Lղ-������Ϟ5}�� P.��F(*)
�l7<B�:n=KQ=B�z#61'y%�!�aW��Ub�H\ۤ���C�GW.i�zܔc�Fj��a-�9^��$�e٨ ���w]��ϧ֗PP6���P3��Wu�/C��n��6��;��f�4�~�>���Ao�!/MZ0�= �4=T�X����[=�j���
!O�ڥo�BM�'���DQ�:���XW}�*�H�a��6:��VAᒶ>�m�	�9r(7��dk=]��&�)�h}�Gܝu��5=�e3�+���*7ͥ�z(�����3'P0���Y����+JG�=ɚ�gį1�[FR�Jj�WRL�~Aį�Ӥ3�;q�O�w�Ƞh�\:1v��_?� 7���s'�s��(�n8p^��~L	�� ��م�p!��������ҳ��B�W�8�v��VhDw@���Soi!���[Wn���)�m��:6%E�&�x|�}��[Gup��Z �~�J����VR7��YP��1�j�E��>L��*n�WővZ�$���g��n(�pwk�yc�֜�ү\���I���@DU6��ClFQ�9�k��e�P�����c��1#'�dU����}���ܪ�D�[_��]
C�̩�����Ӌ2a���8Ƴ1I��<g��Y�l�ǡ��OZҤBէqn�ICN��X���H����8��I$b]3]��N�X��)+hGY�hZ�p��Y�to���I�����9�/.K|v�O����%Ԝ��Y6>�{ΟNo�5�P|����m�pӤ7 �8#-���o�Z��@�cYT��{�x�V\�D�o6�K��P�CY6�Ƅ�ԝ���ϣz~^;$���V���})h��v���_vg�Xt^�g���ϖ����z�C��C0�[��d\�r(o��}PaS�2�H��3�����_e�]Hn�W�4by&�/%�4�C�����l��ʽ����u�7�mæ7����j:a �&4/��P�%g
��wѯ�&����*��2�Ri"������Pn����,������|�xѠ���5�*	T6�����k����=�{�J��,�uj�w��ފ�\c"�o�CR�5��˭5�S��:G��a��H��6��ё�e�G��0�"U�wꑌ�I�J�y�y��i���/��	����q4�6)�~�;T*��2T�!��D���S|.�[�a��^Q�۠T��y诧SD;<qtո�B���ٴY���@C#J�0�/~�GdL�G���qjO��O��VtO:���Fk�-���]o�b��RMϚLu8��f�W�N�38]��^F��0���H}�E����q��5�T+_��5^�%��)[��}8�WmiXլ��%	�\�Z��;�2<j�T�;aK2��ɚNr���֔�8�#�/��*?��t"j�a�=�V����u�K����X��@b�>N��(�x��i&��]�E߫�"�+���MD��-ơh�/����J�8�K�u��z�
��n��}���i+c��|��������Y�TK���;|��n����R�$��r������_�{k�v���O�T�{�H�I��P߫�G6��d��
0/�Ɖ�i�9F�i2�*��Ӛ�?}'�=B[J#���./׆N;����T���l4e�ƌsr��Rw�[������0�KG�Uy��5��0���p����q���O��Ux��}C�|�ު�\L|;��~��#��;�3AM���y1����7����h�us�D�*w��4C!�:9�����݉��C�VkY�.r49�L��H���Sٜ3����O��Ur���v/�_^�p���p�<em<~ҩi�@�������&�qT��m�*Ҳ��"B������*{sS^�*SW�p�����*�bAy�`��w�ƿ�*|�*D~���M�Hv�J�y:��4�w�=O��1/�1c���N���1hٶ�ji�oC�ّ5W�۲�8�X���o$WO=�zq4�T��#J��dak_ /$v�b:��u�w�^�g�}�mG>�%�ڧ���V�K7C�ES�WDg�F���j Z��
���Kl����!Ejw�U��t�/�?���$%�x�jb��	B�N�Ts�e��w1��*���7�N �x}�F[~ws(����ċa��U� ���#9y/A>�J�w�+2�G?�7�w7�eH��ߓ۟�u��4m؆4�'nD�$8^�]:��
I�kaי�������s;\���yw�@O+��XJV�5�,��Zt!x���+�k�O�i���?^? jBm�2�6��4/�8�=9-��p�Z�(iZyy�َ �$�+2��v�,̈��0Y�^���Q]�  ��<��}`�f�K�Rۦ��QHxv�$��¹�HS��t�h�U�KV�6T6�^��d�^C�$q��^��ZNT��
N�AB6�d�Ni��~������+h$�����0+�YC�tw�8�m�f��o(=݌b�6���Y�,d�
��£�˅��h+oBj�����9�*?�.�@��CB&4�3{�oN��>$���z�_І�;r�E���fs�c��� �$j���;]E)wԸ��k�>>����G	a�(?C�,<{B� �:���)J�H^)��b��P���W*����%��o?��4_�ހ���9:~k*L�;:��0�_�}Z�	j<� �N�A*�Ԃe��y�@�}����_�Z�=��B#��P]��	M<���8��Rm�t	��{����sM�+_��؈@gA^t-�f���F*�4!H���#�~�}`�J5w͐2����� ��Z�*�I�a�0�;��^��[g޻N��lY�9���wǗCӼHd�\�AR2�X"'����F�����>��!�x����T!��@(�\���{�5�ٍn���Li�/o Ii]*��"��$�n��w�,	I�Z�&��e2oeC�|{��C�U�u��j�j\�a������J2i�R6;��XQ���X3�И�v��D���w� ��B�
 ����+gy��	��o�8��K5�W�1��a�o�2����&�O]zi8�VOQI���Y6!i/��y^�+b�oǲ42�d��An�(�$��HW�
)��.c�ލ�a��/�t��l�ɃK���Y"GK�ݵ	w�r��uǀ��u�7}�$;�C�=���pU��N�P1�o�.���8����<�xS�>�/����]u1��������	6�Z4߅��1�.�?u��<,`M_d��ڥБ��	 ڟ�n�U�~ťD�9-຿h�L���=|�-(� ����ϼ ;�g���3��~��*S����@&�T���J�;уm;\"@�~�@ �/��yT�{���E�&/Ӹx���E���sW�j�5��ϧ�i�V��Ւ��ё��kA����{N9�0�,�J�����*޴�9�X���E)��\��v Rw�=*�H,�Z3rx��|�G������d�O�
���Ҙ�t�X�'�^�G1
�e�|D��*Zwԅ͚��M�\��^�B�oqcǶ&z(��X�И#��m�C ���Κ*�N9����)5�a�M�;{X�S��Uv���L�����9ji"\C�6���;8�G_n��3ˮ����%щ��o~��j|�N4���/�5V��%f���~((�r��eSj2P�������P�|��E�(~M��5n)�V�w��+��3�� �Z�^3��	��JO���l�ؾk�ZSh,vS�#1�Qv��k,�L�,}�nz��)Hy|У}������N�Y�P�)�������>�g��9`�A'Oww�%n��;�G����sw2Ü�=�u��H����F �ڕ�|�VkeB\���V#�(�Y�o�٤(U���2�<�`~jw������tUͰ&67��	�����t���G#;L`rǼ���t�iQ1�Uz9��.�^���GE$C��%�^�Xݗ����XH�zA'5rZ~J�S��H�÷g��*���E�h,h��r�7QM}�"";���H�X���|;�l���wH��ዋ�r���V^jo�ҳ,bɵ��?W;f����v�r�����jO�̉��e/;�����G��8"%96F����#�E��mcY�]v�߅Cݮ�i����3�B9���"�m�C�f	8�<�vw3��+?�=҅$���r��\�'�l���,�ޕݼ���._�'�g�T2��v�v�%��$�a��e���!uY2��>~%�F������W7F���֫�0�&MSͿ6���D�.�k�dF���U^�jS�/RQ �t�*_��0����P�4 s?���z�f��$���t�������#����;��=\�{M���*x� �GG8\g��T���$ObG,5�~�!��8/�M�ScQF!Y ?ʗ
�r�����z*f���ZG�~ҷ����<l2�Ngp�"�P.Wn��xF��gd:�B�ko^C{��B.��j�T��+����*pJ�ű���y+v)]��L!�胀�{005�n}x�0�yH{W����<83C��}�|����%�B��oy �}��$E6 �qM7�����h�%�s�M5���v�O�8I��[ڀp?\�����]��	eҭD��ɒxJR:�~Ҭ���h/zZ�=I:�k�Ȗ���+�������OsmNd;�i�{a�2[��upo��b�(���˯k]FU�U5e�7��j�S����z�o~i�
��7j��cm�ZGjxVI)2~�xn����&�u�H�lL���;�ZC�+���x���WF�xB
}���Rv���D.�ܝRdK�%PiRk7bT�͇�ķ5�����^��C@�R�uxėx��H�9�H����S5�*�����T�=Y�d/���A�:野�Q
�|W�U��Ex�B���d�κD�G�Բr�	s0������'A9�5��r
]��3��hVʜ1��\p���gV���ϳ
F|b���5��w����m�|��GJ ۴����J"���R*��;�.*ӣ�G� �=QV)J�R�?�gho#�>�vu��_ ��zΖؓ�>��=U�E�����0�g�V�O�&��>��
Kv�7)�T��%K�^!FЖڴ�GLĞ��p\��)�)�����Q���	s�� p�ёШ뷀��ώ�:�I�3}b:�oyL|��|���	���)Ů��S�?���#q�!��.#�E�����=����'�����4�Y��LOa;��)�_эV�;����ɓ�G�+y�y�ey���/�T�k�ϰ���W��_���:ܓI��,t-������1{&�6��&9�#���0�����:(�0�������`A6ł�_vD� �GX��U,��&u)���	��,H,�+��7<0�)s�y�%A'�hE���OG`�YK��߰�rc�,k�1lwU���7���t�h��q#���K[��7��5)��eHk	�%}8a�K�� ��P�)�%��Z��w-킥���񈞜�6�!�=��2�U�[s�$R��}4�(�K���Y����P�����m�����ܪT��,z$ˣ���w�L�_��>=��O�|��ӈo��������e��|֡f�u�"�l�#��gͨ���|�|ў���#�UTƒ=
�|�-ݏ�U@����P�*x[z�A0�w)������-�{4"p�g=�-/<M����
r��z����
��P�M2y'&�O�����$�y�C���@�@`Өԅ	���Km_�s�;��i�F(oF�:�2h2�d�Z0Rf
�ሪ,�x�\���1p(����%��=�]Ŕe>CV/�����f¨"���U�Y�s�ۣ�7�t�	e�#P�-�NQ��&�r�ؠ�˯(�#5��ϲ">�&�?�i�����Q�v7pG�M�r�8�8CJK�C΍aI&RyUX�����+ʹ>}s�����R�U�C����<$�8z��پ�&vCe�ΞR?�`/o_%�oTq"�s_ �U��"6��B.�k��y��:�=9�����$Voˍ���<�{��oM�� v0WG�yo=ףX|K�� XfL��et�v;�87K�g�r��g}���&��5�G�bE��	E�	><�Z��	S\�h����ӹ�������N�iE6��.;�,��������� �b;6�\��P� ��(�D5H�{5�!A)��)j9_xfg����KXHײ:!��(����u��"�+��zv)Mg8�A��`��#�����D���P3M������v�#��r���\�~Ӈ.�N+��C��TzjyD\�����/�Y��w�Ř���H�ޝ5pT:X0�GML=U�į6 � ��g����Y�9g��H��MV�Uh¬u�̃*l>�ڃ�/��(�^6�?�El�VE�q|�31�@�t9!�0+{@��Ԧi%��ۍ"��$8��%T���T��Fj���cMݡ��D�Sf�����Ѿ�51{�@��=A��i<�=���3��X���X���N�<u��m�H$��m�E[����y�"-y-`f���}GV��m����E�?��V6;�sW4�1���S!���U���0N��\j����yh
��Q��+�����s����4��G��NkT�!���n錛���Y�B~~��b�4}��u�ڨ*b�}g[v��3x�u6���45}���)-R��L]��y5�2���Plb��x�!�X.Un�Ý�^�-|i��*�W������*D>�B�%9�-hŰ^C��
j��!��)���C�����Ƕ+�я�����w���5{LaJb&#�Ł��=p+�Y3R�z Ή���A���=moM���`��ķ��[^Ǩ��YH\U�&����U�,,� �#飚%���wI^6�J]��p�0�l0�(O��������w�H����
;�8p�ߍg���ʙ���(	x�;3�zɑ-��.���6A�bG�67�U��U����'���œ�hS�Î�ac>��7����`�(����w傇'>-���EO}�%:��D:�[v�
�¥_��IԂ@|�X��I�?7?V\��;Kh��6?uap��<�^���qyם���/9ߪ�)��y��<�?�g���l������C1��dk��ّb֑�.���J��Dh��j�h�{���E:��i���Л���w����E=e�n���	a���	���������}@����?������S�J��0̾m���M��&�B� ��%uf�\Ew��P�8��H��� �=��1�F%<��NO���h���*����0-���׭�Osh�"�ه�VYli� ��7���?]��r��w���,	B-~�o�~�2����oYCJ���E�c�C[��'��r����4��E��0�>��{؜O����(RU���4�Ӆs6�w�)�G���)��7уklsO��8�C::#����2PId�J�x,���m/ ���)���S��Q����� ����Qt,��{{��/�q}�7�N�go��{Y�&\�I�^]F�)���rǿ�F3���|�مxV� ����wܙ�b2�{���S�����4R�Z�J~Q{��
Y};T�*�-^��_|�.�4V2l�̉m7���B�_�G�K�Y>(/fT�3:�(�-++�+U�d`����ف�}+P��uĢQ\�Zѵ���	�� �!#�bh"q����&�[��U��&?�a
�z��[��H[e+I����6n�7�=FY�A�}Up6�3.�>�e��ܣCIX���(��ڗm#�F��V���VR�[/�^�4�S�+�T9ϑ�E%z��.����0�P���GՕ�@���ϊ{ylɜf6t�iɎ,~��t������/�ٓ��(��l��1LvP�����oF���y3�u5n�N�jl��a�'B�P�@D�2-���h���\���FpҐX̏�^��m��V7F���#�x���*�����m.�\gz���o��F?�'LU����Z_\���\n�V�����Lt
l�d������ٶP������'V�Y� wk��oYg���ƛ�����աƃ�j�CF�ͺ Dj�=ұ
�N�2U'�uQ��R̀�~����{�*����&�K�����_���4�����p��^/�'�<y!�+�Z��~5�'6ۦE���}�Wz��{\p�
��'�b����F~�U;ܖ\����HY�͙�U��o2��٤Ը�r���'�\>cR��ʊ�X(���%�u�N�����*��1f�MP=�v��E/}�]6D�w�$�R:�����=�[L��0Ɠ}�-C+Br5���=�̮�H��j2�>�ĠN!����2��1��o��+��aР]I�O@9�>��O�d���F�d��֌j�~��Ey؃_�A�b-��Rz�Uy���6�T�c1wa��]�&���I���zld`]NG��.��޾���B�WO�������[�b���ɈzC{��8���_-/�9JW��
�!魙�`<rtG�M��N
�a ���}f
��|�o6���t�*��mOF!B?��i��-�0�ZSjXK`Ι�	�"�F4;��?��h�t}+��	�x�7��o"�屟
���������U�L�4foe%ZF~]�pꀓ���8\xd��gSs2C�Sc��a��D`���V�z�Z݇f��D����ڽ�Fc|6T��3�3�����r��MF��p���O�n��Qr����X�uݲ.ڽ�F����g����\��.�Ra�}Sc��Yt(�ִҝ.
Ζo�J�ȇ4��d�v�@�rjt�L�]��yr�wl��:�`"�g�����}�:$�e3�W�qV
gx�h�mۣ�~��ׄ!���F�	�/i^ME�!h{�>5f�Xֿ��)�Sm�|�חh���oWډA�O���E�a�oY��P��Br��`�M⌯e���	.�%�y��˴WM��4���Kk���JDg;����ٶ����jQ�CW�+]��9m��/ܧ��a&o�E��4+D����+[Cˏg"B���-4����j4_R`v_#����N7�\�l��xp��ݡ�I-����,�����\YJčv�L�ԩ�h�Ͷ�.fYM�F��jt�U࿓Ȗ�����3;�� �?4�(����+�����z�<'���N���͡F�nܼ	� K�I�C�Y��_��xH�׷�1D٦�
-�^ǆ�e�P@t������H�ԉ���3@����*�_M�Y�Td��pg�.�P�u�?ZU��Q�dx���,�W�2&J�h�q��;�O�e�W�݄��v@��Pf���
�4��%�@��s�;�ezYx�~�S�3O ̰��	\	v-�[+=T��m����3 S��G�kh���Y0{h�<a��w��7{�`yƲR�D����1���O4��,sg[��ڡ�:�V6�-�!�d�FQ.B�@I�V.���й1{��*f%q�n2�g��<�������0mz ���t Yɻ"����h��?~�c�^�@���΅�d�sR� �^Y�!����B}�ހUDϰӢ��/�)��)��u��lw�%�<������R7�-M�	����xJ�m�P"�n�j�)G�y u,Q�9�ʄetx�Ϻs�>[ơj��%���v�B��^��Q����P5��J�F�Ѣ���u���Lm���?���e@�}ᎏ ��U/�4����%X7'E"�\^�3MM��Q`�ll�9�!T�-^Ok�PI\ku?�X��9u5�mF`.ꛮ�Z3SW|��&�l!B3��W���Su�o�B��+�6��Y#{�b��*���g�B���"��G&T��O���BQȀ�$�@�IZKCg�pA����7掗���6�R�t�1�F�hg+��|���x����5_�.�K8Lg9���W�K��얩��љ �ջkO3�DZ���@0~�F`�[�c����X����9m<ji� �\ ���u�>� �		�	.�cv�`���.:���"	�{`{ �{��JD��`�ч����^A뇟��Z6���AQ�DC6�i�����*܆Ϙ�^�
�T�S���\	�n����#ߊt֟�F��Ѝ�Jnp��H�&�^�I����D3�No ��]��$yC5����,!����;��
R�7���Twg�:z�aR͕�5)Q�Sh��n4۝�7���S[ލ����qE��s;i���0��+y�5VP57ܣ$��mY_EW������>K����5t�|Qa3�{ݘ$sI Y��v��}G3u#��Ty-=�s��j�u�ϒ5+`�t�j=t�6<Vu8���(I�x�<�lԭs5��&4@��ʼe�(�L��ZjW��v�Aik��e�O�Ψ���͊�;���$}�@
���巯�6p4�6����e���Z	W��n�P��70m�^`�������qL��g\��B��;�Ԧ���ŝv�n_|��L}�	�ja"D��U�:<���FF_�j*� ����Z6��e����I��渡��^��=ц���x�ˣ�{����{Ŝ�RS�X[]�K���,E����^�z�jo�����^;���V���/o착�Ů�~!��-��W�ύ��z痴�J�9W��Xq�j�g R��թ�04������{,~F�Tc�g7�5ǹ|0!@�@�slI��eה�X�r3��S���4λ�6�V4���U}8�t�]LS��%�^0�6�h��E��i$�n��{�W�  oۉFM�HSb���<�������c�p���4y#�\D�웵�n��Z== \�j���$��p+��͈e$H��{�d�L����+}�|Y.���͕ON�#�oXeǰ��t5ȼ/ק�ԬV��:m�gŌ�Rh��r�+7}�O���+&"�b��6��np�:�Ay�t���@�=_�
��ր�/��&atÇ�o���/�/�Pf�M��0bU� �6�Q�/������o�����Pغ�ܨ�6��MK0v�M��Tu�uq�_c�M ������uFz��"2���~(撍1����YHB.2���|�T�ű[h����q��:�%�3�+������MMs������Wq��Z�n��Q�h�p��P>h�AL�ۓCA�� K��O�f�KGR����Ql�;���N�r�/�]K�=���9�H����_��7ґm�2/~\L	��
�ׄ�^(��W�
���	�h�ѻ���9�yXکPNR��G��������k�Y ��y����R�͈�
^���R�Ĺ�K�mq�u�낖d�&>u��%��J��W��2}��r�|����2D�϶�#��8��>�t$�N���*�U��g�tY_ӥ��*Z�=�&֏|���Pq�C��	��Ü{����P��	թ���Hq�u�ߣ�Jjp��~I�&4%ߏ��O;_`vX�������q�[�}�G�KԺE�D�?���I#�g
nY9̻Ze��o�-��������s�Ucz�c�Ge6r���_ޕ���R#������!X�/f�P�g�Y��	d>���ٝ���
�F㤯�L�,Q�lꕸ�<����IK���K����b���w�	�p��2��e���t4�&���{�q�O�� an�M��Q;,K����ܦ�9����'���� (�����0Nm)>�}��.� { �T6����r��0�f7&�O0�����;�R7��_��I�?x���Y��Ca�4Segw*�X���;ρ���X��?�|l�(�H��ʤ�;�:>Ӂ��ɰ�!���mQ
8I���d��kX�`��v��(�|�������Ť(� ���f�6A�� S��ol�bQ�c�n(��;�|������v��Y7w�jAm�Zjc�#���޶����<J>3%�k������i� �9"Vt�}5��-6=���wHP��,j�Y�DG�eZ�̖��w�
�Mo����`Iٹ #�����AN���Z��k�Aۖ����wXK��K�Z˨���k��|/�A�֥}=9�B�jK@#��!�a[;�Z^���!�C�+��G�U��?3�J	z��sGa��8�M�cKo�[���/�C�����k�G��G3x�fe���%�@�����HlW?P)��u�k���a����A�frD2�m�U4��� M☜�.{HhG4��\�Ѹ���q��n�AB���o�ZN�7�9��X������S�I>��U�cg�8**���u<� X��K�g
����N8��^n�����H���Vy�J�JbQ�-|wf[��5��A΄y�GV8����2�y��~SG$����Y(�}�D�A���ɮ����1kN���sX��]hj�ܮ�R�5$��$� �����n>��r�p�O^�G�X��N�>���rfz���Po���5h��_2�e���(}�ώ�c�D�̖��x����~i���.������i��?(���+�Z�?��r෿E���}�֑�7��[O�Ҷ�1���@��_Zu��y�R�-ox��?&���}C`0���__qnq�`�m��w�F� 3�r([���H˱����l��&� ��_�2[�����{�WH���k��>�f��_���L�+B�u� �օ^/���Y��/��X����j���O����S�����P�8ξ�ɚ{K��p��z�k��)���"�vʱ���=��2�y����lhR)��4��9,E�We���t���:o�CV�Wk X��F��(ˎ8C���͙#���9*b��j�-]�_Y�4�PS5Ԝ$s3��y?���ET�)��2,��~�{NH聧�;��>W�^Yl�a�*W&�����ܣr����^�E���!�f$a
:h��6�[Bt�V����%�c�׆[�uZe��-� lYY��k9���۲p��)��I�4���NAt�4J����N˵~�5t�y �Q�.�*��� �۷��/���7���ʿ딻:�tM�����n�G��5Lًa�j�����9ϗJ����#��>u�tsN{�V9�ʋ=��E+',#����|f(�(�59�,]z��D��!m�߃��h7�����F<��7�9�cu;���3=5�cʘ�o
�~<u/�M��R.�U�D�bQ
�*#��8uj���f���UŊ���1[��y�Aebr�]�W����'��"�}�$h�����K�6�Bc7<�v����8�~��a�Ze�t#�1���/�!����� 3�*�jg�*�<dk{ū|ƨ&|^ u���-����$X%G⼵]�|�.q|>a+j|������nz���La�"-��^�|�:�g�E%�g�ĊO5<��j�X;h[�ҿ��:���+���T-t�[�E,M�;"h.��7���ip���2�C�\"|PC������X����rx�X����\q6vo� (�:cʸ��!�X�:!a��ؙ7R��t2�`��T� ��_ =��{�T93���3�m�z�22�n&&�?��_����&A ��\��Y�#�h��_G�l����8�V���	�n�û��C�N����c�mr^J�L��G&�E�˺�.A����N�z�L�H*����C�@Ϙ���<�)�3�Cvk�v�/$�FN�=n	�82�_陧І��0{L)��{�\t�:c��gv�_ɢU���@�mW��3���an��g���w��78 K����8f����\���Tw��6�%+>[�K���ɧ;pJ�&9z��{��Ӆ�M<��_�J��kG�̽��!��g�m.+sy?��&!&I�Ǖd$ƃ�Rj��*�����!�~z��]Y�E<�K^b�]�������b�v�ʈ��u�E�|g���n׽�? jь�H����~~tHE�r��`5��pؘR�;���2.�ʼA�;�rj�� �4�]qw-W{�Qs���c�L[�����{`i�ӥгg�Ֆe��ຌ��g��Q��*��[����f�Z�_{Gz(��8_�d�|	���-4ۚw��W6,�\ɹc�?��`UO^��	��r���k�.bDr�.�py�=��HB�BV������F8T)���$�C,1�������/Q	�BwK�z(k��ʟ����@]s���v��_h�m�X\-�ɾ���`��z_Y�#�y�\��-@��Ak�J�JO9�d�Lْ��uCSú�^#���=]�uiK�Uͬ
����#�#M�Xl��ʿ0��b~��F�l�X q�{Jq��#f">R� -�C�$�Sh:s�+{"@hKP.���+��#��������_�\�Պ�L�Y�ss�1ı�V/����xm����(������Cze:�b�\�`̞Y��3�T��u������w��b��
@pقք�:JБO�Agp���rb����h��B����7�� *P��9�Ӳq�/
�EzUm�x�`��]�v�C�G�f�S��@Oc�skg�.C��y�b����� �,G*�#��jzli�"���AC�/�PhW�n����_��[�OAV�;G�H�5��q}�Du�3�q`e���[־�;����^��H_����9��g,,��v�"x�������6cN��]p:|FZ�|lN!_>�5�Ό�@t|�E)�ѷ	kA�Sen;'k6V� ,��s��[��U�!�f#�@��C��j8+�$@}}�OL��{]�e����^�� ֱ��)� �s�t�1�+�n).�:n�(`��*��_��$:4�����S{|����̄���j� L�ӏnPb��f#�/�rk��CL��m�G�o�1��˼�����z
£ғpy��i�]�D�]�Y:��S͚�B�����QCd���T�3<tcM�n�qk��[�r`��qI{���� �R[U�\�J��H�f���
lV����#��V�̹Koe1lQ���7�5�10�%�I�_�$!�b'o�X��t�X�py� :K
R�);#Ib�:.H9ͽQ���*c�X�=�Tr_]���%Y�2D��d�o���D��NA*k{{1p�)lA���#a�N	�~��4@
NZ���O�	�l��@5ܹ+K�y��$�y�Z14�~�6ֺ������q烆����J�s�l7@�΍ج����;B��j&�?Tu�����FI۲<�7ķ���YeGq|�X�?|�n����K�����Z�Q��Y+�o��y�� �5Tb��?� B�t�� ��wפ�)ys:{#�IH_Z�}k$���w�!K�Z�΀���Q��w�Ek�̾u0C��5��m,�Ġ?���D,q��
V��D��s��C�;pd�'k�1�#�d�� a1V�f�>�lш����x�'��M�+�m��K�U�抈�����d����\.H��o!�e��/��)��gılu���y�+7ͭ�,p!����[�P;�o\M�i85G8'G��}�%OA��I�Z���K��\���UѼs����|��K?��w��׾��B����4�jbcߗ�s��!��kC���-�k���
���i��0��49y�t�G�&T����RF��?/kn(ĞU+���.�[N�>���i�
%�ۆ��vXo4��3�t_ �'�dnn�F��';��; �fPmt�-}F��(�@��D��7��;l����X3K�4�s�
L��%POW�7sH#�|�[ҀO�� ����V�ό3�
z���2ϲԶ쟚y�'ل���GJ����3���]kY����"M�����+�cڑc'؂��0m�d�n�d�ȷ�'�]ck.�"��2.u���9ң��~�u��YaC�"�/�d@�G._2�+�H��.��;
��ĔE)��O9> ��6���-���?�l�衬a@� $��A>���5���4C��4�8��-U�|[����`lm��� _v��?���e�9�;���nN� p�M(��QG\^�X��Z�0���$���
_�J��������^dS����`�܏����˼�Y�	z洦�QGQ�/��7(�y1�����e.���L*<ѻ{�*��sd��fW�#����|7��杰�j\�2-B��u�Jj�s`�Bc��q�]��9�����ű���ͳ�D;eg�x�8Aש��*\�F����D)���:����K���e��r��RU���_V2�Ji�o4���]´��(�;CXӪ�j9�ŦG�O��W��[�����2�`�e�&��#�bW��&>E.�D�P{�;��Y7�7���e��c��YQP	ay����ij�{�I�v�Q��8���hA����O�jYڐ��x�u�3����%��z1��+;V/�V6�l�� ��ꞥ��IΓ�5W~P=v�s��l���|���D�Dw�R��i���5s4[s�#g!ׁ*4�\
�ՏdN�'_�F�;��τ�J5�[���)~a\C�o$/`f���,찍؅8`I[ ~ ;h����J�Q6�L��QTx�Ҳ�>�f�<��.{���!��@$�'Kg@}�y� =n`��	EV�Q��몵!n����F���㑋�����\�6�P>9�W�G���t��7�-�a��k�m�M*LuY�$�ˢɿMu���̬�,�^q{�5���V���|���	�Y�P�C���s����ފ� �-m�f���>|!�;R�7�9� er3+�<5VC�~�*�p�uf�J4���_��,�ca� j�`��U�8������j������(��~���NPК:B���hl��lZ3(�(�i�? _�Z�@k9m�a��̌f@v bb���8x�'OD�%�RxW���ݩ�a:�X��iG�evM硟�,9��t����vw�,�ilȾl�O�^��Q<�wZA�V�(C�(t��s�+��7X�)�%w Ԋ�4Yh#�,-3ӆ�ߍ[o�|�o~+�K�L`�o ��h�i%���=@�m��F&[� [�,G�q�gv��ם	�v�V��y�~N���� v~%l��t������'Ӿ��q�4�a��
N󴖙��+����+~�[m&��s��0��n_�gŁ�S�0��nJ�6b�T��X�yѡ=nR�_�w���b��ݼ��x��y��4thq��'���D.n����"&S,Jgǆ��ڢ�����v��ĖM�pd�~�:>��Vڊ֣l��y?����C Qb�/-��v\,��Oc�� ��������8�y/�>AX� -�G�6�ad�or�$FP���O<.���_{r6%��ۮd��"c\��[|o��t�������^�ް~V��� `5�م�~�Xa<��RS�����	�;���!ڭ_7��Sڣ*��R���u����V5��"�L�D*�j�(��VǐCp=^EGr��ec9��)�! ��vbzW�֐�Z]U>m� K�g��S�Ԃf�O/��oi���vy0��f#����?S��~R�`��v�18a������7�eۿI���ژ�2��9S'�;QJ4x��x�@Z�6 �X�f��pb�0+a���i�f$$�� �}j���H�0
f��[b~����Ŗq`���_��.�%�޲�ȅ���><H:���W���Ƣ6�3Kjӵ���ʩ�I�4׌騬�'��aPn�������Q�
�1�l�M�?�K9 ���v}���ڂ��b��M��57r���z�!����u'�����2$����^��#�^.?��I��V%%�Z7�b�0 �e��������~��#gn��İ������4����aP�X��1�'��)���bp�pA){L��I�,�2`N������(��0e[�|�\�@`�� ��d�[����?��&�`v�B%Z��ZəX{p�^Mx�yX!(��&�
v�xI����8�/��;��ȷ����?�~�X�ϊ6��L��3��ڳPPߙ&�y���A�z4i����$��-�Dy�KB�Q���v�ow�E����,f?�b:J�ǽ⓱����;E/:8z
0Ӵ��Վ�%��`tLw���OW&�cmx\A<J���֣%�I-�u�K�s.<�Qm]=R,��U���~'ÿ�m�N�ŵ�R��� ���n��vh��0.-��>��cL�_I0��|��i�'U�r�K؁�oT�l�[s)�?O�0Y͘��'�5fU��0�p��� G���Սm/XRMn����HaB'$=l� �'������%+�jAAhл��ɧؙ�\>����n�b�ՂS��^�U�+��5ML��KSU���f���M��3�_!��S�x�����$�� �"$1Ffl���#�)�G��22θL�X��H-��={���+�y��<���G � ��f�	~�.�#N�����H�5�e�ڧ:Dp:}@�ζ���EV�j�7I	�����J��%"_����m��cL��@K��wF�/����Wl��E��G1#̠����&��j�5X6�M����]Zs�;vp*+���:�o͉Kƿ �ZE"+�:����ޫse�"Wn��|~��BU�uh�/�����9�.vH^r@�G���)�Ԏ��VAl��n�oT��5�`(�2�R@��`��"�jyJ?��R�e/��MӺ�NV}M�ʘ�1�7͙��M�=�$�C3�%N�}U��5��B��zٲs�)�Hs_��+8�F��w�9IM�#a��g55��Q����2S｡n�V�_V6,����[	��=2��,�Qt巺�x�n������'���'z����!���sT'p�r�%cr~C}��Q�I��c�S��Sw�ɲ!qB���tp5�-�[f��߷J��ݼr����IA����1�(�;���tC���/��%=ݻ�6�k�SI�g��@Kq�͎9�V�"F�z��-Ղ�S�Ť� YJ� T{fe�`�+�p�P\��K�Vc�L�4o��� � �i�x����D��i���1h'L��O�5$�%X�oq%��_�d��\���4�S+���r�J�L~*�ؙ�"n\W�j�xc$^]���l��'��do�N^'k��ϰg?P$,	���>������sk�MD�x�8�Q���0��x8Č�s�QE�n#g5�ۯ\M� ��Lg����e �O� ^q�1���w��i��	�k�����(Rx�g��uQ���D�#���vk/��d9`,����u��Mڏ� *����O�(A\C�UX��w�1�|�jH4kf��V �JA�
�"4CM ���ʍ�>�{�1���O���9o7�M`n$��U�b��L-.��_��,��aI�^�f��9��+�n�R\�")Ƶz�/��>�-�sY�ܟЖ��u�\c_�d
�@0/��6��Ѽ�@*;�ڇ0I �Xg��������%7�^�/FgRߜ2�
@Y8*���`�2�J
L=u��EJ�m"mZ�Du�z&cx[�	���U�޿3�=����4���/����R�D_��~ڳ��O��-V�9��S��F�Y�ܣkﵨ��EtD)��d'\�$��t�!�����(�7 ��.B�A�0E��$��v�\M�c������S���1�K�������m�a���D���������نwv��~��V�9���u�H�~��g�H�O
��R�`�'�{j���:�ay��-�^ē�� �J�n�]E�ݻ��t����܏�A�1��;
ո3�(���n��"[��
�6i��C�m��Q�v���/��u�L1���m|���'��#���C��͟�M��i�|��톱L�ᑽ�ed�B���`J���x2��N*���Q���J4j:�O�S���H��0;�?N>�O�����Y��
���$���d\�-�E*�� #�a��b-��]*"�]�j�4�_�C:-)z�T��<��v'{]��=���WI�/^���z��(U�^��?fB;��F=�w���g�U�裻(��oMڒ%��ų|+0�W�zvѹq���d�؄~(�"a�jT:�����a
�V�)_^`��;6yU�
���m�J����+�cB�3��zԂ�iK�?�:��?�ӎ�F�ܾ�|��3ĳ׍ua���E��|ߗߥ�+�ˑ�^��Q}_�/ϗ��ު��
�� ga�}��3��g<�DP�8-@L�?n�z*�}��s�f�S�N����4�a)۳�|�(����_)�����c�1�_��/a39��EV*�v�%�f�}6@�1m1 �7�X��LyIqvW�*�h	����ߟ�� Գ����[�ɚ'v���0�ni�V1r�w��	j�b��^���$�����#A�
|��ht��'W�D�H�yi)�(PR:M�A^�	�ȟ(O5���QhηҨ��_Q7f4A�>�z�-�Hǒ&�K��5�_f�e�#-�e���;�փb�\/Q�.W4���˪�CM��Ŷ�8��ż�^)Ұ����"|�RS�T`���e����py)b�d����1/�IC�u�`�<mVڸ�Q��(��c�PT�P{DP�G�x�ԋ�*�¹��7>l�H/����s��̷��PB�5>(�*�i�d�y�ȐCZ����T���pr8������J����L�#/��e�*I�~ǈ����R�ް�]M[�C�!��e9��g����ȁ�:uԄb`ٻ�u��n��Z����x�x��/6\�(72'k���l��Aoz�l�l4�v/S�@*/=�A�8������_�U���\�y.Gʚ�!�b�UM-wb�_��B �P)N�,N%֘d�J�t-����&V�囓;�%���I �)��X�{I��c������3>��q�z��V��t�����|R�G��,�:=�uЉ;T�aT���<�Ƨ��|q��ׅ;pm��'SO/�z���e��%mUP]D[�6w������b����Yޏ3vD�[ڋ�� �5��^���j�Ӽm �Q1��fyfW6��C>S��Q�N��.�L�qjCe��R�:���|�����0
N���>@t�믪�67�_G�X�Y���V�(o6Gd�:��y�����Q��;a��v�j�d�ֲCD���j
v驷L( ;zVLj����8p��`�vR�2�V=�P�Gp�}� ��Dݐ_/d����)��t:�t��� F)�P�V��m�����b�� ƒ���Qe��@;Fv?��9�� TO�Lf	��1��������)
|�{�͋d�u�m�4N!5.�L��sz�7O*S{(l~6r5���6��X���^�V��67�)x�: �D0X�`�J��i��9 n�L�X�a��OՆ��e����J��\�|�:S������w��}p�@�r�ؕ��c�֑|Z�����7��n�	����Ny^���쩥�"��J%Ñ���&@�A�!�GU	�ah[�!X�_��}���qI��]J�ܮ�V集��3�T�/����7i���u闱�׬����QK�����"�ƋtQ���MV��
b���Y$��<=���Kt�i�`#aW��Q���3s���~�vJ�Z�{��]���RG��Θ��.�/Pq��V�>�##�a�>?k���QǑ�2�[U��W�D�a�&�����'�F��M^���#{'Sf	w_�?@�-���&��.�,��Ə��1y7M���7M1el��H36�݉y�kO/�ڴ��.��&��,Nܥ�Bϻ��Y��
�6���oIej� ^u3���`�$�0X��CT,�ˇW����~[lS���ˮ��en���tp�4�u� Z��`ɠ��B�N�$9�iJ����v���;t�װA�01r�����Wӛ�&0�=��=P���S��ګ�p���%�FZ�~F.;M!q�j��O��/�9,;��#��rg��[!�_@�+��1��o����¯��sG��G����:�=P۸l����W�E�`|�jb3���'�t9��;�|�LWjd�o�_��a�y�-W6}J��׉��b9
���d��|��X54N,�^m+�D�"�s;i��(Hp�i��c`/jĶ���e�f�x�d� er�@to�����p�[o�smI��@�֫C������)��>
�l�'����A����.ԟ���F�c��Nd�p�F�� �w�%���ܨǹ�N�\]�pJ��F���{zI���9hC$'����Q�y��l��	���	�4���\Z6�7�ӯ2۲��[$�aQr|/H��F��e�c���50��41�|E1w�@���� yI�5�~��Ƒ�`I4���V���eKB�M��0���К�����U��"l<���r���£��wĺE�ʹa�_vM�[]�  U�;����i���U]}e�U`����4#�{C��=�"�C��ǒ�v�OI�	���;��#��Xʝ�<1���S��v���������%�X#�T�r2���
���F�z�tӊF�ϳ`�\�k0�N���J�+��v�������$2�������a���S@Ha��(��>j�"� l��w4�ս��V��с�����mН�2���Gҝ�^-��O����@f��+B�<-�z�2wX�Y!��D ,�׃�)0�����2FX�Pak:�X���P!�%�)��5ZQxTG��e��Y�xZQ]j�m(|Y������=c�Z�R�t��w�sP)�6��l�QFiT��i�aJ鮰�)��"ⰴ�:�:bd�;��J�� ڵ!-��w�d��v�-�� ���W�����C���z��������Pr�[�[I�z�_�S�#1�0M�\?ш����g�� �ճ�	J�&(����u�V���<�q:�383p�w��($ �bE%�Q�����pn��.2�+�OO���2�^ֱ���:���?�P�\b���o��ʻ��E�,�HL�0[F��������瓌E]����	�v���՞V������2I�ھ����4c�
�tm���gR�}1�u`�����9��/߼�p��jQQʹ�j���wuޥ���Gn��t>�>�����O�:����v�WeL�<p5���cBfAh�ee��mq�jM͆h���5v#�Rv}g8���0��cn���q��^*p����X����ӵ�ko�Pc��oN�=u����G��ϧ[r�=�,����'�"\�`��{�I��#dd/��5��*'"��GQ��XQN*O3����A�`�}-�H3k'�i�5�Q�pW�Yޏ,r�  �G�u�QB�B �\���-�!�e��4�,��f#��M�q�[�*l1�����k��8��2>9. ��&�O�B\��?;����I�xS���w��W�,��w��*}�a:w�%f�7�q��C���p��>�͛
l%�n"����pI^X����=p�?����TZ�V ���%Q�k���l�B�"|r�m�Q)�&3<s��?�������R�zc�P	J���-?��z�B���C�9�V6ڌ^�0+�S��p��jq|(�
���CՎ�!��ףepF�ٞm��唑L�tJO,�׍hg�PI�~�v�A�Z����ش���=5�Kݶ�ݣ��3��j����~�.�3�{�����kt������h�bet�`ع�99w=��9P��e� z�]U�ڗ����i@�3�~��X�����F|, B&9������a�Z�*v:H`K�����MQ���<\�m�0��1=�%����g���lG��A�����l��	貑U�h!�U¾�����+�eC�'	ґd]��F.��m�>5Iٖ}��ur�EaƉ���ք ͫ�h�ψKOZX���X��v�����tŗ���2[U��@�EP!���(.>���w�c�ӱj``Q�a�u�O�s�溦ǖ����+�mo�-�H3�8�����b�����Gpʣ�'�3�.5�D�H��Sߟ�X��G�H�~�X�Aҭ����'�xJ��J�����tY�9�)�}�m���ټ	p�mïda�î�ѽ�a0��grb�xUrxo���X_�V
�2(=��_o[�3�JN��$���w�*��;��&X�h�ϫ��=��QH�9@�u���pي�C�Uj�,��v	��b������I�#�̄u�\��ђ�_Y3;E��M��u*�O�����Pf&#�ƾ���u���[K��ۉ"S��to7�'�[��G�'� �P�šP�>�r�X����_����vی��a��ϥ
wTC����܃=�C��uI@���052t�`5�����-���K���p���g2�N�}]����u쌉�xdXI�����SH�'�2�uh�#/4�/&
��[�Ƣ���O'���'��4����w�f4�����3��x�1O�R�b���Q�hƘ�4��ɕ�Q��]�Ѭ^!":��
x�;�MT\]�AD�@�V6�􈡄��M�M=�J�UaG�)��~|� ������݅�  Cz�`�AMg��Ŧ��g��(�����#vq�1�%S�_� �2�`a�?�lk��[�Q;
����8��xpz*�q�ruC�,��`�)J�<���p���oO
.�dz�5���/K�xX/r�~@w'��Σ1eLՇ��K��T����Ȁ��<������|ne�7���1�K u�X�Rԧ!�2��6eX�ͷ8p�#�')FF��ť�t���\"�;�׶x7�����Ĳ��i��3u���o9K֚)]onx��9��#�dӨ^���V�/�b5�w����q�u��P�o"-�p�a���[E�<���t�f(�������-ٿ�$n�CK�J$?�������"8lxN֬_2��dc܄Oz���wp�{�n�-P���Ї@��?b�:��q����¨G������J�U$��‌���a�(��vVY4H�pJ�Ipo���o���?��;�L��p���A�;�<|�ܟ~�xz�d�=`򼾠���gb��w=���������g�����XA��ݹDе�V��S:�����J�f�љ��L�BYz��-��1�}��/��v�x� \[�i5����Ƕ�m�?]mb���fN����jM�K�t�i�{��_<�NLy� �9�6�=yQ�.;�;�>tyVK�Hc� V���j�<��0�x��8��.:�)�K�EÞ�I겾�BO�,�)N����/�������<��꧍sp�YX����l���)D._	�qs��W5Ɓ��FFg0��b��v�/�4�~n� 6e"�N�"����2�,�2�(S��pF��m	�]�$t�k�@�#o���,�A�vKcb��\l[��@2��*q,9�"pCN�����ٷ�vO��0����ë�˸9r�����hK� ���j���fM�S��o��G��E��f)��R�뜖�@�� �3~�P5DC$�c��j��[�F��k�T�x��afݔ�U�l/���E�Q�����)&���u� .���2n)��G�Ĩ'����3��	����f���#|���N�KPCc�0�?�`'����5�O�A��7�1㲍���ƢV��x��M*�T�����E�H�ky���"� ^H�$�m��r�:���WyߣKN���Q�pԶ��������h���wN�TH"�4����p��&Cm�0����jk��bj1�����er[yA�.�d��e�é��g��#�C6	<�tc?@�����;zdY���Hyp�=O�'�`#���z&*DOT�|�Y�����)�C�����"�W��dׂ�&�D��M�m:�XyZ���J]D&��y��k���܀C8��~��y3@������-�`�R��<-��^ܸ	��	�x{�-��5��2��<�ף���� �!���U�W��@��lB/�,�N��?I>*�n��b�j�����[_���;7�,[��X1W1���EKw�<G0Z�����Z��$��3��@v���I����D]���~�Z����(F����?�ʷx_Խ�GT�7�ǰs�r�����&G���	T�����<�����&��]¢�6>��1�G��	���
�9�GZ x�+��t�^,C� �W���\-h);��j��yT`�
������sָ	�g�2��m�\��m7�D��8�Ȱ���̧}�{�����X�x���y#~��/�XB��*�ȝ���̓}%O��[��pd�C8�� F��,�{�TkԢq�|��r���+ ;�2�M{Ƽ^LLj��]��J5	XS����ugUPS�߿�������)�csH�����r �2��CT��HRZ�-�1o��)i���+� I�}���k�������Ƶ��=�M�>[G�"VH���d��vQ�3�+ă%�.�Nk�C�ւ
��Dr�1a�>���ՐMI^�{m�dy���m����)_w�Y�4�W%V��� x�ÊE��-ئ��y��t�`ht>!|aψ�>"<l�̢�����k2/�j=2DN|��������L\� �H�>څ*��dz� �(�שo�'�O���#��B�N�l��z�B�]��Ogq�@?2�:\U��w♺hX~ ���5o����[�:x�Ts����-��h��RC-L�c�W���J����`�e�I�4K��ͷS����H���77;���,K��@���~���Aܙ�8i�J�DG��L��/^� u�C�F�Ņ�)�b��Jڏ��^Z
V�GU�+��l��^����ƶ?0�t((Π\%6p������T��D�Z�{Ʉ��B8L�������J~G�}���+}��J��.��&��a�{��}�/�Ik�~����#A�1�>? �?�!�0�Z�v;�!�!��=���ޚ�K������ѭ�KFR\j����b���}��o�6Y&�� �4n,�����wM-8����n�W�g�BHG"�I�ٜϢ�n֢y1�A��ĖZ��d~��<�4� ��Қ��&��6����u��:/7~�b:����W3�ʀ�O�	$W�y"t�lˍ@�gB�շ/ N�% �t;tR�BL ΝC)�ӑJ�U�'#7��e �����/]'�Ķ����p9�)J�־�XOm?~����ֹ�����y&8Z�,bϯ��K��O�pB!&դ�¾}7���d��+���U�#�w_��V��m	@X�g�B�q	|��|��p��ƪS��*_��<*/����!�3/�s�Xu����fH0{I��"tq3%�3.|%���|*�@�F����l(�hX�Lu�\�.�\���-8F8��8�YU:{�?�ɞK/��*3x�Cyc��ϜԒ8K-�8���=�����j���EB/��~�Мꃃ��Ǵ?AטXD�~����R���{��㯵l� ���X-�8�[*!����OLO8���g�&N{�O�����鼸�� ؂GE5
z��(tRr�u� �@�Fk�C�X�k��[�������	Q=y_�֫�Vb>��^ڈⶊ�L���a��nL�i"/7V!q�P_k�IR}�e�#�����e�xA��`�1� �U��O�k�i�[M��m� ���� �r~?��/ "��U&��wVJ�R���̺j��X����ĳ�ޒ�(�'V_c�m�9�u��JEL��s@�y\?�Y]��J�A��L2l:V��zb������z�������pY��mj�<�(o@C	���8�,���٫�}��L����Q*F|�m2���|�cF_CB_V�7'��sE�y{��0��c{�M��:M�8�ZS����߼9o��
��[q\f%`-韻���4���)�
$=��C� �0::euN�ZL6�������3i�/� ��N�C�yB�V�q*�������7�����������c�D?�N!�ay�	Wt{����j�Ng�E�Ò��]k�1��P���=�d�.��zͷw������s����)���L�,Яe���/�Z���f9��Dٝ�\��=�TX�%�ɬ_c)�V�<Ǉ��)�u��Eh���e	qV��
K��gd�y$"�i���MuYޮ,�0�P
t�7N����68����c��րe}��FW���vz�E��I7�X�)�U_��^b����k�Q���J��Yަ�c�o��葱�����k�Rp��O�h�)PnQu�k��h�&a9����gX��;l����ȷ�����Ř�q눰јR���D*v�l�sf_h8��'l�qb���������]�$����wĠkQ8{� �k��9�2q��8������R۶�f��PTG:�o~'Y��a�@��!�r���0��]x���%���Zji��TFvM�W3�3�J�%�ɇxMy K��ۜ��aC�̬}�T�?��5�X�L[h,��(�ٔK�8�^[�\�h���O�'v@$��ta��A�&h���#t�|mܨ��w��Ll/��m-��&�F����I�Q�ɤj�o�|H����Ň�(���0���$_ܻ8�xNf����K2Ae߅Q���Ɋ�������U������ř�ԟW�F�}�}3�/�́A��3���*Or�=X�uT��\�]�}3w�ϛJc:��Eu��CP��Kj2��+���ѢB����JY��T<K/�m3��ky���T������oG��yk�w��d�������Jd�)�����`����q�(32Pzڍ{��2!�<�'�Ʌ(�`�m�h�$�v([7P�X�T;����,ui&8}ą�6:̷�"�N����bi�0�QxRN�p�������(D��)�r��i���4a+)��<P'in�h�=
A��,u��O�|��i>E��*²*���Bt��[���O_N�M\�Ȟ�jI՘$��6ͩm{֧Q�
�����e��Ib!&6���o>�Gˡv��e�Z�%�<��*��aL�TV��v�X&���3C��1Ლ�А�ɦ~�"?������/�z��ϻTG��#�3L?<�^f��[����4m��n�+U���Y8����KB��N�;�`��?�/����x�z�A(GZ{�����l��Ŭ�s	�X<FkPʬ=�����k��F���j�Q�Ѓk�;ſ�v;d?s��\�A%���-��c�[�;��7�D��?6��Q�3K�+��]1߉��v1�<T
v�}i����H�%E���4bz/��h�Q1N�����ܴ3+ۋX��d`�R���:�H��+��h�U��F��4�g^�����nk�����*H|�^DC)>�I�_��M�L�^d���ژ����ϲ�鷺�N? +>Rdߓu���{U���q0�(�{ ڥ���2e�mgZ�x=�ގp�ܞ��C�[�R2���|�k�@ �j|���$1h��q�a�t�ґ���y$�Kz�7�� Z@`�g���[t��I3���q����\���G�қ�
�N�92s�*����:��@%�)������4�
Ft�mV�R��n�>�a�m6JZxC`���+�P��h�OEsg���rm9T�	�H�E@�Ҷjx������-�����|^B,1���=ns�Sž������z���nk`���)��<N1m�ľ�����<&[���^׶5ew���X����7{��s�:��A��	���)>���������!uN�uZx�����6��L�Kbhb��%��B�>�Wju�0�O����K�FnssqT�m����DD3��V���Q~��ٜT�7�A
9X�פ�%�� �lyx��o�"b��]�Y����3���c���`��|8%��[W�h�*���N��)g-�W��,��_җ�/$��<T�'�j%��{�M����~42r"�Ҹ'87�����7�`�o�ƹ�����޽�>�S��N
�����t��K����Qgn��v�!�W�>��?�M�9�1ȟ ����DN�1�|z��g��{+��7�X3�� �)��e����҆Zg�+>vV�^y��i�S�|V���|d��K�F�7��d�
i'et�����6���o�v5�7����)ZA+ �������>fꫧ��W�=��"m#(�Af�[��N�sq�
o��|x	�権��n`��䈢��B����m�ܻB�%�{ƴ�F@��R���:<�m�tp�|�IjW]�">��%K����a5�8E��ӝ5�� M��(�Q�,j���.L���0��==Es0����$�/�nE�$U[P��N�W�F��߼���z ���J��H��&�ZB��yil��\��j�� ݹܱ>>�M�:����랑�5�4�}� V\��������P��б!��z���`��Ý�����n����J%�!�ʞ�r76w�qsUq��d���Ig�(����5���:��낍�Y���kF
��b ��ľH,"�zN�am�|�Q��АV�c�(�3w�A��,����� ��!"��=��l㚙)�U*���\�� �8�����ia��%�kT��|}�>#�d^���D����.c�>vV�n�zq(��sw�Sp;>MP�C���jn�J+U���)�շZ��(�6�*�b�lD#2�-�7����3�4���Uo1S�F�p�6־��2��ud�ч�������~ٻ�H'^rԌ��5�klmD�aӘx�ɨޤ1����@���j��(��Ec�?� ��,nL�kg/\�P��oĻ�G!�o�`J �|b�M���6�k�&YB�;͟���ܢ�{g�k;&;�J�B)�.#XƩ��w�	�MΪ�@���2��-Ŷ�?�{���EgG_��v<�"�jY�'���T���`t���%4N��ƴ��ENt0Ηo�2�_g�B�µ�xP�4 ��s�P�0�p���\$�GcH3��I���M��E5.~DVӶa��x�}k��lփSj�0��❏?2~�s�� ��3,-��߃�>�~��`���Z�.:����L��w�I��$�:�5>ؾ�n����cƱ�ն��AD��;�o#��}cO�4��!�.����ڊn�#��xVt���0����n!u.k�T^��˰��؟�p����i`/����;n7�В1��)S��H=���V!���r��٣	���!�D��
�D��Ԣ!\?G��]F�=v��j��`�@c%c�X}#lՠ���+͒m5���
E++	u)��u�~l��.�a!	�5���L[*���6	B&-��X�+����(�f8w�P�B��X�7H�a'���"i4�2]�ON�J�=,	@8���?�y	���:c��Ώ��-A�tO�[!G�ZSP�h4;��HD����!U*�Џ]j��yQ/T��|�Q��@*y~=�I�ϱ�mI�P�P��ۺrF\��5�!��¿y������Ҽ��0�s����{�FPm8����ƶ�&���)+.��
�	�o�ٶs1�F�DFH+���mL�3�<�S]��O6u�d(mf@�~q�&	���]E��$�o�	n��U\h�;�q�}�k�/�j��!e1,�������X�}u
�[#���5�xđ?;&��he�9D�<,�jo��J�����8~"s�\�]��vR���=\U����ێ��]�j{�g��oT��/4i|��)���~�)!��V����S`TY-�<�d@�'����0Z��:����A}��9e{�9��H]y+/#@q�����7�G�{�C�At�oD�D���]�e�P�����92�E��71*���Y��b���N ����=T���PT���K�v"��h4�M�D��Z��m�!��ܵN�����M.����I�������G�q/�=�t�{�'&����|6%���89�P�Չ������%��*#�����^�h�	��q�j�E"�֋:P��Pp��1���^�nX�_���;���ڶ��Gr�������%���� f��Ϛ�#�C��P~�~va*`��A��{:H<܉-�ǘSp�'wt�:I�*[ɓ�_x�ܲt1��ǩ� �d.1�!��\�"�,��v8<��q���mo�ăK"4�5��/U�
f�r�*5ЧBw���⣃ub�вzE��Q��F
3��73��q���-����5���bP>�.�O'��mϓ���:��<ʕ/�yd]���.��d�$��C[n+ߜ��tA����H%��~��	��z�0��}���j4H�q�טӪ�� �LS����'\ �w��x�\W��tn�x�Z+T�(8����	�!T����&�[QΎ��"-��� ���P�  ���Kj���X(������1���!P�^�QM`/�+�vjI)qj�/P�p*���xw��䙺}H{J򊵌�R�5Y�h�:�����Np�'X3%���f���u`@V='��Dt
t�!���:�N[u]��`ݜ=Ң������y�ywԸmF�E}[{��&���W�B0�!�fj�0}.�j���(`(�j%D9���¤�1t�Ǜ�uj2(P�s2�^�����	u���.�F ��D>���q
?���U����S��\(n<@�k�<��g����]�XE���|"��� ���j7������T&��9�
\!��D,ug���A1�X�KvGz��!H㕚 ���<^6����l9N��ky���	!Y#��:>�ЁKV>��E�1�w�*S���(e5�z0Ar�O�Y�����j��
;f�i���^�~�Nɹ��2���둱��TEa��3��S)�^�,�Y�F���Ɵ1���R_��v'ao#�!e5���ח��:�&M\���|ss��g����DY������'�Qn/*���ЗV�]G�����W(T��j����J���NiWj�-�2�]�@,����}��Zn�_c�U��mRT�@{Q��������LfV�:F�Q*��r�4|WA�:�g��0a�c~6<�k�G� ��N��n�_�W`��p+f�6�Bl���l�~X���zE{������U!3����f�o���|��m�:�{�������j��� �Q��	/ڟ�$9�u~0iI�����fh�<�����o���շ�$�|$m/]�XN��/-�@���S���2������I��r���lz�f��@f�� �� ���4�v�u!6���ajn�(�$uS�b�1�k�rnt������/YQ��� hŜ����#�X``�\���c�N��{��Ø'���?n�"(+k��:+0�G�Pi�G�ۊN��B�@�f6��r�A�nzB���K|!��RPN���Ž��D�zI�q�ks]�����sg��1�!�� u��2�����=��p30�ie�<�HS��r�3�nf� ���n�E��<��R��Y,1����p�]x���Q4���R�j�,ք+�uRw���b��-�G��T>}����$������q�����'�;z�F�U<�������MC7@�n61|\�O��C� �6�2�ѧ�br�����q��M��|�1���`7Ph��س�`�t(�EΛ���rxᏬ�_{����K��3r"�M�eh:6�f�zi�p�Ya"aeӔ,�@��<���6�j=>��RC���'1�1 LT��,7��(/kQ?&�G{&̐��'i Q%S|~�!>I�Q���!V<y#��4&�+-Cyۤ��j(�ql_8�o�[i�-cT�ʃ
��xЄ(q��>挴q�����f�jU����ͫmOp�튌8N������^5�Aq�/<
�Kw�{�إн+5CO���#Djg��֬�t��-���9�ȼ�Ф���l]��F7YGJ�8)Y��]K�r2w�f,pj�l.Y�֮f�U�&9O}SD�<7��8�䠾6�����<��(5ul�%rCy�d��3Ⱦ���5&bu��_��Ta������l_����,#�h�tB��'&�Ǒ}G�	�q"�|�{�S��m�>�"z4W��t�QJ%�Ѥg�t
�ש3X�S���8�q ^9�����cjeY~,����C�l�A�^� uuo��0���4�x�9^k��� �v@��$��n,`p5Թ�gu7�i�UC͛9�C4~��چ"�|�K�=�g�hr�]��i@l:_p���:��ʞ�i�!����//=qx$j�Ċ�Ukx�T��Q��֧'����s�Lڹ�r��i|#G3��P�����+��Ύ�X�P��2U���h���u��^Vr���t�ƒ���AL��j2QU�߫.��U8L2YMR� =�jd}���r�v����H�e�}�>��Yy�";d�M���ڊ��~'n��Y?��²�9Pb?$�x��y��_���wq�|1u
��g
;�j�G��n�����W�Q�p~Ȳ��q�g5z��n0�G M����,��EB���.kY�X��!��HX!�qx~��!��Y`���Z�daq��G��l�7g���1����Qa��
K�*}��k� <������2�-x.�Og7b@���Q�%��������\X۔9G��K
������D/�;�s�ʳ"�s�ù"��;K] J�]ݝ]�U\�P�ŉr��*�}��I�J�F�B97UcCqF�����ԯ��1?��W$t6{�ޗ���Q��E=��q���Pr=b�Bv��*��G|:�k�v���bS��t��aQ^��f���B�T&WǍ�|���Kb>�e�HB��$Y�� ��>L&��2 ��{�}�p�f��CQ�rS�dߓ#�d�	���^%�g�z��[��3���������:7��VƔ��������=��d��5�M�y_���l��	)�0x�Mu��WB���T@X��}3˟���,�m�k��7��*�\�r�X6엍l@���O����CQ�5����]�*Ȟ� ,��u���RM=w���)�x>��i����8u�	y�.ȕJ�Wfؚ�S��EƁ4fdh>�!��n�U)z��[ �7�G]�qF?���v�ϮDx'��Yr>-Ȏv1(NZ"T�{���ߥiّ���,�S���z��5/9��q�ء2�u{͖T�I�#�N4����r�?>�Y�4 YHq�x��y�
��)e�u���.j�F��%iH��{����������,Mщ뛝xh��EZ�'�t�1㻇���"֡(T[b�x�.N��~����)I+�LOGu��ϏR�T[�M@��>B�rs�i�u��#�h�6�_Ӝ��<��͸f��\�>Yѡ��i*6|��*�����~;X����2���}���b�O�i�\jm+6Nܵ+n���Yl�gz�|qD��e�Ij�����=-B@��]oW�2��Q�{V#_Q���6>[,�e賝�`N��^5�38�Jt�{��R'��G��޾���].��!y���g��.ɾ3�<`)O���u�w&�:�ڹr.�$H��!M���*�$�� ����I����i�&y��,|wt��bƏ<��5[��l1I-�`�$,�N��`���Pl�}PG����Üg'�K2��=����l}fw���x"��V	�	Ҙ�����GV[�r���ؐDT+ �6f>�d
H�F2�Go��Y��~mɶ��<-G�)[��6{N�1n�j�����&�yZ�-�oM���ս�	;��c���L��ʤ_��(�
یЄ�r�A�?੖���AS�)4���!���@�.�b���ûqS�Q?�������R���'P|��ˁQ�<��
3{ǂ�ӿ�909�stF�F�k��G:����F �*�;�M�6�9��"r�}R����g�aY�S^'8����^@���w�K��H��@FN!���񁱈�����Rk�i�2X���f�6_�zʪw�Q^@d�3��զ��M���Oӵ����8��饰�J���q����\G��.��(ɖ�l�e��Ņc�,Ż����7����n�j��g1�3��wGf͜���չ�+�)�z�|n��!��u�&�����h�K1�%nz?�"��&��6�s'�n^a-��SИd�aϪ�R��4�m�,�i?|LW-d��rB)l��^P��&�R~(����b�Ψ�y6
��X�8*��(� ,�\ >�b߼�+{ۇ)Ҁ�\��GFI��BOc����1����&�
��K�HC�/a����۬/|ʹ�$K����G��X4�7�Fɣ�ƥ|�^b}�^�@��#��Ŵ&�-�"�Aj���VT���cuI��n�}�"C,zw,7���-M��`�[%3OY_����D���p吽�=vK�aS6X� ��F�M���e���� Ǟ�e�=
9t�1�� �}|wo��u������UD��/.(ܪ+���Sh
�0ͤ�f@�����s���xz~�7�1x}�p�6�J���LB��ks��D�TdI��̈́��2%B��c�'�}9Զ�Eu6��!��S�oC�\�I<S� ��ʎ� ���KdU�>���.w����/;p� �m��Q�Z���[~Mv��Uc��';u����Z�e�ܕ$�{����>�W��� 	�֠�C��h�q�>�[��*�B���N�
�������G�	4�F���0�@��ɌZ&ԋ!�;f��9�(�^I����:wD٪�]��_�a"՝&�< I�T{D���������b����B`M�=�L��K���j�\4�:7Ԝ�Kc�������&�~N"������!讖"	Z�xO��ܫb��l�9��fϏd��.�BCg�>w!�`�R�OϑO�YȈ!�j���H�,U�����e,e�'SѢ��-M��:<�}�`X�.��J϶�"|����$�_��n���N�m�(��X�j|�E៩ޡB
����S��C���o9��T�:�0�;�3��'�&Q�S�~F���i�z�O����/�@^/mh��	~���$���i�{Eh2^���ąlA(�R�Ɩ�?�u�&Y�������-@��}OLQ����4|�_��,�?X(��"�ӟ�R���.rƧF�ת��aӚ��EC�<U5�y,C�<���e������
�^�Ҩ��k_X��cR���$�������:�v+۶���KI�|�������Z����Sl�}O�~6և�.h ����H8�i�Y�E+&��r�ʋ���1]�c���`��HY��6����;�JV�:��,ɡ&�h��Z��㾱�s#�9��M23��歏Pb���J^w��,��Z�����ZЎ%���:ÿ'͚�p��Ɓ��x1<թ����!��,*a�R�b�f�.gq�!a�ϽHāp�
�_�"2~/�@�v0u,�o�m��QE:���e��|����Q����ϡ�82�v�R��U�����[tU�
�Ρ�fO��#�#ɫ7}(G0��A�Z��+wb����
�v=�@nLw���pT�dH�\V$�J^jp�-�������^v��ղNmZ�(ߌ��f�.T g���YK��r��n��I��^	
�+7����x8���J����� $�%\�&Ji��бX$��S�E8åG�lm�1�?�L�NL���z�w�Z޻��0>�l���ë�6�F��r4���y��ͣwsg��Ќ2B�k;�R����\Yzv_h����qsJ3�9�F\� p��@����˯��0�p�P��u�������o��O��<t�i�'x��Gd�2do\�%G���%���v��!	̱����i�P/��Rh�6m�`�#mۑav��'���o[~*2^��Sr� ���=��쎫J?�P��8G��.�c�z��<�6�3g�`���@����̢!�^ѽ�e�������b�'��_��@��N� 8�(�3�v^>Qw���c⍸
kpQtx�f��ƥ�J�Q�N�����w�/&�O<ȱ�L�
���IN���V�Q'�*����������V���*o��Ϥ���Z-���.YIA7��ۏ�ʷ�7Q��h��0T��V��n�����52��Y9�j���rf��q7�j䏈z��9nhQ%>g���;� ��Ne���z�zH�u^We�h~�(���B�GG���Z��lz�웨(�ӝ�i�<B}�,�_�rYaTR<}�X�_	@��ֵNC'�:�O*�l�$���8�`-癫�<+đ.��1&+:���C,�%�t���&v�Lp���;2����@y�ϊ9������r@*ٚ��<�x�Dz5w�N�#�>]���`5�*����㎣�	S�{Ks�\rn�-!n�C7ۨ�N>� U���b��>Țl?���f�y*x^spf��ɾu�����y�ʢ��5B�X��Aq���c�-_��K�K����Q�2�M�e6I5��%(]�����[�Ɇ���<�*�I�䄈Up�-1�7�ݦ -�Bb1���Q>oa��S�?��C�Ot�W��O��a<��Q�y��CM�m�}��=R^ G�d}��dN�2�ہ��2]nV����Qq��4 �AT����6�Na�&{������! ������|nߤ���:9��80����ڠ:z*��i)��`n~i�\�*�Pp�����z�:� �N��=n�N?#����JMV�S-�s$�	>!|/��ւ%j��� �����~�|��<ފf��0��'4�����x��w|�X
��Ш���}�q���=Iq����_�.߯[�Sm�[�J]���2�pAB=}��*Y�T�t��лT�TiY�Y�������]�������>�GyI^h �o�`M,����T�Z��>���藥���c�R�2�E����, ����1;���������J�ԬA�s2r&)���G;)��o�\n�����%��R�?^&������o��ʉ�	�e���eg �֥SLۄ��8e���Y%ppE����桺�شW\rb������
��EB��\{�3�oK�p��ͬi���,��R��W+;�����]E�/�Iߚ�,a{��	�vI7�(� �r���"��p�$>(n Ǐ�L���l�i�u�L�Aɠ��W��W�W�)k��?�}�}\��;�)���������ܑ���"e��g�o����:j~ɒ,�/���V�Ԝ�#�E�ƪv���*�0���f&���9i�Tu��G�D�^�<T́1܅
�?߆$�"4��b�QY�DO<G�Wmَ��!_�3W��P�B�s�OyR�P�bF�x��أ��si�rs����c篑US:Z:���ҪO0�wm�|���#fN���:r�P�̜qT Q�Px���w�k!��>
@�H��o���h�����$�ϥΉ�Mܔ\ɛ��zfôP<�k	�-�(�2 քs�o��7���h�� ũ�Z�Etg�Ѣ"�`@Nt��uōͫs|���H�bOI��|ܞ�� ��p-�R^�-$R?Fc���iữ�IS]���ؚ��po�V:�B;i>0�A�Q���YN]n�+�5��UO1���T���6!�'�u-���ݩP�8�"�Z��	3�z��G��G/G�dq�a4��ȳ��s��6����LU�I0X��P)*ME��d�yz\�ac!�#k��K��n�¾4�kF��Ϡ�B��b����D��2���G{)g��AF�Mڭc���t��H�75�� 55hIE���D� Q|j�͚�we-1O��'�,4�2����M?,�A��@��Ǘ�����N�5�^���3�՜$���[�Y�eM�vf����Z����}�GHj��m�i�K����pз�����|�٘e�)�~�|8�)3��1�lژi��I���'~_4Xx#�#�=3�-U�T,��B���4���k�xx�M�F8�_��ʦ����|~�3�-МD���T��\��h�UX|XF �񀖐�[m�|�+�kA��w��������'x��sg0�x\��/,�ӵ��)G��ޏ��s0�����!�Ft�~KH��g&��̆��ܚ�E��x�����ޔX���
wY5���HO M�=E�,E���Z�r����� �y�ɤ�¬�!�#��s�s��A�o��D�>�J�����P�Q_K�#g���9�Q�2��K���;��T�\f%�~���;���m�VBT��!�ثCF"$�⠐}ڢ(���+7"���6'ۻ�s��IL��uHC�̏�Z�n�	D���(֠�"��1娏��).��f��΍�[9
	b�d[�M�4�Ն ���j�Bn��Wx#�$��U�T�3F��p!�߬��98i$�P�0$��
����0�Ғv*�M�X���	{v��3�Kn"��U�!pY^���$��ڤ&�2n�n�!ᗓ��a�ɹ������[���1�Kw�_��r*k��|�՚Xk�2�� M5Y�S�6�y�B�nulV���i��L	��g)�Kn0�B��)�+i���DQ�3o�L�6�5�.����t �&��RQ���Ћ�z�䖭�dW���gl��
W����,©zD�޵<�[��f8��\��QwN֝�B�W����&qAqMY]#W�,VmS��������'���88F̈����-o�i�O٪�hW~d��?��ҁ�V5��	�����_XO���>�jg��m!`� s��s~4L��Kg���u=�*�]/�4�۶���#��������W����q�2��|UG��V��U�vT����X�+W<�1��Q��.[d����[��4R,C��S��[���� �/��'L�X̌nzTA}&G?�	aѷ���ݤ���p�}C@�w��@5{�1	��g�*QE�]���$W}����N�Ԏ�F<��Ɗ����͛O���3�ǖ#�����:a��RL	�ltw��(8���ԛN�Y�`� �d�xepZs]L�]��~8Y��2tw��У��T��I�e6�C�\Aw��t1���Cw@Ŵ��G�@&L%�S^,v]G	��P��4j���uኛ�{mB�s��Z>����d�s^��������M1�<�J8dx�U��k��}��*�q�*��X }ԗ��-ٖ�,�x nc����Zn���	j�����4A;K(2�sK���o�_H�Y;s/qN�.�Q[!J�{�u����\ s��OԬ�����%�r_�4�k�/�\��ۇ���̥���`�**�R��S�é>Q�h�ok	�vJ���B�p��|&o�b��i��eZ)bY�w��M���Yэ^	97!��$gV�F}����Eʍb3r��6� 	��hG�>��b��g���C�,J�6~Gs����fsK���E����uˋƎW�#bN����G����B�Y%�I���sN(�Ou����[��h��J��o���C�T����{�8U�j���W�����ȣ���]�9���4.�$^�.W�*0��B�{z�FFI�ǧf�4���2���y��M�P��3�'�S��\��"�6���.B�[��ΧP��a�.i��_�b��Jq�F��*���M�G��~D�	����Ulu����z�}i&8�d�!V�ˍ�bua�c��B�`����Y�X8*��c��B��	ܣ��U����y�%0�E=ο�h�U�Fnmƾ\��kxD%�����(�s����-[H`��B<�{,�g��,��!���%���:�6�heՈ|.�tN�[��X�k���D~]�z$�L��O���\?$iI<'t��+c����߱�{a�d�vT���0<��# 4�"�=�'״\���0r�?�̀�e�]E��ՌxK�U�m)�O:h��}��3�%'Z�t���'��e�YF�]!��C̫��w��ya�ʄ��K���X}��1��qFW�_[C �.���]���qE����O�Ӥ�j{���\��`{�kk�I��fGk놼$ڄ�!���c Bs�~�T�+6K�`=��6Hg���Q%bue���6D��;$��i���b�E����k3� :��S� ����H��<�¨�tʩ�_`�1g�&��/S6/��F�YN�к'ף�\�>�*9R���߭���Z�D�7{��xE7u��$�r�z�N�g�S|F)�j�;RuZ�B�ߚ�d�K�ʩk������#�[�`	yn>#d�Yi�~]�(/Bހƨ,1��=�M�4���������~Ǒ�A{��O_��eρ�~��Is6L _��v}�d�$��ˋ��:^s�b���43�G�V�K ���U���Z�d�Z��װ�m���xy,�h�l	����I�j R6���������C�Z����bF�j}�:x�/�D�ͨ�?��B�0�uAq?>)�Hxo�2��"��T��?TP�$MCХ«�~�����?����~v��I=33c���o�:�I4N�_���g62f>؆J;��π��-�)����.l�`u��BlOz=��c��B��_�����rP��3�C���(u=+�w���W��$�6[��}\*��x�r��8Ũ��ԇ�:���ZϬ�}	W�~P:�lD��*!�1 	�)vybTK��v��5�D�H�D�Om���轔��8^�mT~B� ;%��n�HoE��r��^�y�p��x�A�:I�� ������Nqu�j/�k�n6�(����~Fk��8�@��,'$#[�J �L�v�[�x�o]�I�E��$��ż�A���pafK'j#�G/���X;� ��>�Ѩ��}�[����ٜosjDo"��8Í~q�p�^�-/�%1Cͅa�*>���B�d���[�o#p���Xf\���AΧ�Y�Hѿc$ Cv'P�T���O��+�\����_	���.C��e�M���r)��.q�i�\��wA�T|�����N��<��M�md���v>)f�!(�J�ূ��o&�dR�JԴ?o8��2��oc�ϩ(k��|�Oi牎��'�y�n�bB��:�=�e!��m�9����!i�7���M5�˧RI��9�ŧW�9xܸ?�O�f�GtV@˩��b����=�j,�מ[t-��Q��J�\_ן��Sh����7����^�f��p.(y<�4x\��nO~������=2W�|ȼ̻�a\��5�l G.߃
�q�Xi����ܹ�������XN'.�Z\Z�<���X�eăJ�/
��}�~	�Q�yc<,�O��IaZ��α��cl����.(^���5xC��ZѴit"8�ܺ�?ҷ�Ŀ�L�U����yiÑ��JG�>�H��ȇ3�ĉ$��M^�E�S i[�����i3�`s�����L���wu��q��6��Fa�����I�^yC�]�+S���)�Ri�@9���@���K�e��:�@���b��c���X�b7';�Af~�QzZ��݈�����������N&[�#��T��$�V�����!����g�h(����0��_���i�����"Pg�h@�K̼!>�&"�)=K��"/Ɉ�ܿ����� ������q�;�y��V�d�u��%�0re��ԈY��
�3��tI�� ��J�&����(N�[�N��5����$>�[i��g,��~*��KHf1l��3��>�?��G�$T�<IÈ1�&�O��\8�.����S�E݄Gs���Y��ם��!(�̥�`��P2�2;�0Eo�v~���#anU�չ�f�Y��	{�E��{��2�u6ކ��	sL'����ߏiu&�/�K���h5���8ܔ =$^��V%�y"��n��̭e����(wx����4s��	W�=_��\{��sv�H�i�7�����#���vY�u�輤V�.��D����)�p���UN?�'d-7O�
G�ώ	P�H|�dʚ����⎉����(zO�%��Y@h��zR�Lyױm����+r%�T��IsuRpQ��4���-�s�$���3h�uk�0M�-�S�F#iQ����'C6�ρ>�	͐|�����~���Q�GG	8C���'5�Dn%�t������y��ğ�*gu�<NU���12�"Cс�\��jj(� �l�w�o�a�~���=���yp�W��H�NC)�;�Fx�� �����Jh�Ǝ ~�G���nדlAlQ�G���8� A�����z$r���ƟK��%A��2T������5WG�yL��*Y���&T�������n$ ��c��3".������۷n����ʴ?���~v�A�
i���N�C�]�em3�G���s}�~_!� ִ�u/�4���6A��T.��\5&a0�������1��v^�5?4���@d_Cxh�Q�R*�0Mi1\��FԮ��$"x��
�����v�h>cx�.)(��B���EW�hۆd,}y{*�T�m,X�s����XQ���r����M�tc���5��m����-iɤ6��#�]Xo.��\�"�Ǉ��ڙ#=*��3`C�v2�U���ꗩ�����KRs���u1�*?UɊ�5�-4�u���l�%]��1	�*yR�q�"wu���u�:�9��m-����)��sT"M��=�Eq���a�^b�v����b9����� 3�SɧUB�P�׷�Ǚoz��=S������o;�I��gFNnM� �j6�O����+ivzF�#֟�E�f�p(n�.F"��@jvu\��t���>�»'x<֪%��)ؙ�u?���d4],<��?B���	A�������Po��2�yWhĻ��7h񓞾9�B�����U��t���;��|2�?L��ly$/�
Gۣ�0�k�,%0�uq��\�&�9R���t3z]4*�o	x���c�l�]�Uu���"�p���[��jk�y�=��*|)��rb�y���>�d�KL\�"&Q5�����8�Wt10� �GDn��̹�>���/n�)�g�t������h\��"�;j��c��@ḻ��N�e>]O)�M�n�9���"��Q��B�Ų�v���딕C��sQl7s��_�O�,^%YR�7$�M.�7Z����0�W�JP���=bI����eⒶ�w���v^��Z	D�'(��c`-�ÿP�R�S����';d_�p(g���Te��������[$��N��w�;���T�N�Zn;8�:��"���9g��сhO�f�3$z����6=�'�a�X��;ŉ'VFBⲪ*09V��J/.���7�Qy�i|�f��#���c�vĜ"�4�#R��W3�'������L����A���QzE*�!�mP�fs,j�!���49��7�$ߞ+����Z��qٱ����b��Ζ��A{*���g��m�t�@m����ë��o���Ҥ�q�Y\�:#�&��(\"�Ykp�m���_�Z�>Z�E�l'c��}?O ��	R��RԼ�ר`�|�}���Q��(��M�U�2���	/��,*���,2����U:{##���B<o��Dk ׎"c���|A�P�-KQET�ݏ|��ض �&�	�X'P�0�9>�����y=`֞�փ[�����|�8Wh������#"i@&����ŏ�H�k�V�u��'�i=�l�UG��^wl�ߧ*l�%"���;O���&\2�H-�}���+�d��Wj:��	 "L8�Ǜ_��HI�+��K�%#{��?汜&Q�"��Y��o�n�*F�� ��Zdy�[�� ���ٍ^��6�<�tވ>���ŝS%ti���V!#ݚm���z!ٕ�Ԟ�	�/�q�L���v�I
�_t�����P�:+�k�^��H���Hr�$���]��MQ���g�$����'��b��/׫R_L�R�ܤ\��έ�H�- gf#��@�\grF�+�(C3K?l��~��Ll����W�a$y2&	!D��c��Vȥ�7��}R��"�s����j���,;�V�򒤊�Om{� bg����2�+k�,�,���{H!�t�k�-ʸ��(�δ}��������Y��a�����z�=�9�)��[#X��QS[V��W������>U���f�kT/�&.�}.]"�
�b)=
�k`����q�ɦz�g���i5�Os�b��ɕ�� ��6z�^%��_%��x�F��a:�,���<�ex���x��^n��r�;U1�ԠϱY��FJ���*�:��u�����qI�����V��~�e߯cOq3�(������[��hu1�7E��MhL+��F`���O
��Q"�����Jz�j�f3��!`�KSi�H����F��#��V��ô�Ǘ��E+�9�`"?��j7W�s��` ��r��\ϹN�[z}��"�څ�K<ք���7^���9�Te'�Obƅ4zfݪT�yf��'������D6 q����b!M9�7�.xK�E��$�_}ْ�|��4�Y閑ÂN˨�Zi-'^5��mC_�~Wi!5P|_���;S�@���:��{9gB'7��<V��W�G@a1elnz;HM���V�r.�(K�磄茈43��.�}׏�>��8R��%���Y�IB�F�`p'�D�F�ֻ>p�����$��H�L�.~�q��z���IKNj�� .s��_vԚQ�v L���~5/��_�~��_�=��c���"
hߟ�j���	�����na��\3�M�AY��߮���� ��������L�
qOu���&�X�x���(��X��9�^���W~'���@M��r�w���ϕ�Ea���F:3������c,o=RN�3���>ay��o7��G���¶�H���H�߿%��a?�����A]MH�,��i&�D��򜵷B_�Y�z�׋R;h��?bŭ�����E��4�&�v��j�$���"����l����B,}1E����1���4%ϊ� �/��)�8�� �M]�a+a�}���i&R�dCR�~萒�Pm	�䉸�Ʌ�xP�,䵸@����"���nm;d�������|L%�	j$0��[5F?Co���,�(	���� H^������^)?��8]��{�-�5��ϗ�>0A��)n��j����*��](
q� ���Մ���i���@�#qH��3��I�UX������w�#0�R��]58�[2f��]�߬�4����3R[�.�vR�x�sU�ɡ`�<�.�jt��|]�����}�}�^v�n��O��z0�5;�uӈK0���k~�.�*y�< ��S�D�t��/�.���][&)�.Sv*��IV��))�(����BC��<�<т��/W��[�t��s�6"�.��>P��Ln��(����[�Y�SV��H��B�Ϊ9��J�	�C��K?V���w6H�ʥ�M�E���bj~���9j ���^���xĘQ@���Lμ^/[A�g����q/�Ni���������%Oeް�x�:˗�5�B��J�}������� ij�ƃ$��'�8���xB���S�Ԫ)�<�B��ym�wOc�k�8�'E1:m�\{I�d!��|��\D� �f�O,�k��t�����˞���\y��Y"&�#{����-��nj}]�M��!�����֕�*�z�$a� 5��@Pd&�� �a�Z������Bmd�lr����	��FZ�e+ 3����fY8,i�g葧�YS�&f�bW��w�;��Vy �(3���#=B@l�Bp��٥�}�g�5�Xˠ!�H�`T�o��s���4
{�ηG�k/E �.���*'�N�
��Fp�_yS.�Z�YKg����w�`�����a3�ʈ�W���
	E���֭x�����u�t��)��mV����J�����ߕ,��t��bhӰ���� r߃.c��+��A������zyC3%������Rƚ.����I�r]k:�?0s����n8��=��=BE��� �?�~��4��@i5���8s���q��A�@ӄ� �bcJ���|J!Д�Q;�����Zva����Z��&�3;)�0��m�����9v��P2�����yW>���ydx�h�V�l�#i-����@)���(|�T-�X �c�,a�=��Je�m��L���0E-���:fZ�''� F0�]:��=ib��®(��/"��l`H.��������s�eA��4k`�e�X�P0P��[�Gd�S���fU�Uɞ�`�}{���`�C��Uο�C^u��%�Y6��!T�Fc�6��3"ԻL���p��u��t��De�7��l)���ӑձ@�SO7'G>2&�t��n�s��C
�_�S5��u�+�N!�AA���10G(�rq�>8`�RNYE d:�����`�B�gM�U�k�s���i�,�e�m)w����o.�v�2�HU��cx�H]ic?&m���8�x��8��6S��jF�����&�_��aΝ�$fx3�ܲ����j_}W)��5�UYTZe�o���K���Ȥ0��3�\�/M�?� �,,��&Ŗ)�4�I�-��[O�_
�krx�֊i��gRG(Õ{~t'Q�8���9�+��ڼ�Bs���W ��(P�v0�l�nx�kS{�I��H��[���AC�a��|�}2ѣ4���f|}�����cK��R��~F�rZ�����W�=����\G���*}��;��u&ѵ��ty�>����@s�P�����+;�>��`�^�]"���9�K.r�Y6[����0������T�|U��:���a�5$L8R�Fϛf�A%?ݘwhn"�JORh����6Dp�����q��Ն�'K�s�ӧ-8�i�+in�A��DI�)�a�1KC!���`>>g2>lZ�<@V*�c���7�e`�ieo��x�m��c#���=7~��Tf|�7�{�E�I
�텯��`�0	®�#��N�<��}��]Dk)Q�B8�m �~HYk1Fz1�ч���SR`#?E����������,�9���	�	pMc�*�W|�����Y.w.S��C�E)_'�t/`Uyy��I���j��"	ئ D���q0�R`�|��R��r���1r5D��^��q3�M2d���E��]���r�),�J��*̉����h�Wm�m`R��$2)-'Fm�Ceg}|>�Q@���<�5�]�z�-�s�����3����7ʝ*��v��K��{�+*KS%�@r`�a;����n\ֽ��o��[&ِ_;����b��z>�d�� X�����%�ޢ��wu	Uַ�AS��Le�k���ѩ��` ��lCO�������O��I��p���a�򓋁2��_��L�����=�W����'	��	��n�=1��ɶ���3�f���2�2����3�%��Bv8O�YW<��Z�7��ơ��Zڳ�0odr����ʊ�p����M/,��K����E13�YBQ����7r�熬Q�dDu����a���6��Tg^nz�����_���*Ds�FЩ]��c/a���W�ᆂ�T8�N+�șL��>t�!�eB,m�K������\B����C�Rס,e/+ߛ�����r�|�'7]���3�Y�i�`'n�
���5,`��8��YX2�T|�1R���F���Q�/�`�f4�7��[L�Lf����Ɗҍ�e������8s��?7�Ct|���秦��ꄥ�8H ��B����jH_[
���QCFL��}��KA^J'o�Oa��(9"@�5ġe9�5/ь-���ȩ!�w�̏Wozx��C#^!��@ūK����(������D"�� �����O����v�tSF�����b؋6�Y4ͥy�c��,��ٸ��N�u:Tfu���9���O�I�Ys��h�>H!�"��<��!��*��B�Z�)�9����	��T����T\�P{�Pj�H,sÂ �Ʋ���4��2�ؗ�J)񬋪n������,-�(����7O=��v����-A 6��=x�/<a{�+LG�����ܸ|NnB�cJK�Dtn���n��s�fN�Y_�K���v5^�����P��|úK�y&y�w< �^����=�sF9�#��JI-��wsIN��;��*������i�	^��� U�Mo������.$f��|��'��#"�������S\��g.���Sxr�+%K�u�(F�B��W��Ku8���o��:I!ٯ>"�QJB�DW���5u�X{G�����x���ɱU��i����>�3M�U+����b�WN�1�7�[�V�R�6�j��o`@�/z��q�_�����5�����Ȧ4��0ة��Ǭ���)i�G�=�8u��T�l
/W�;�J{X��q���(j���bVKI*oM[^ N��,b��1\S���/�p���{�:������_�Q��j[�{�QE�J�� �N~� {׺��*�װIq�Ǳ��,�~���%�WP۠N�b%|1<����/7��v!� �l��M&la��h!�zˡ#%+Jr���m��q�r~8��KDt� ���Lي�%d�$��1���~z��3�n�̉���D��9��>�x�6���P
A<2oB9ﻨȈ	/uJ��iu��M[����R�t�E�7H�0��ʰZ@�������p�s8��y�<3���gq����'lR���:x�O����}�T����OiW?�׾��^�x�c��ĒS��'"3o�ŗ>*�܏M�V��Z�FL\Q$����*���רCT}YrM
�H�6��� K��!���Y�� t���ft�l���(:ʰQ����вdv~���x%JǢZ�Ȣ��s��^_)$�*���5-�<�y٘&�<&�˴�H�T��TO�ptu��F�2���BVk���X��3ag(�D>�N�9��p���lAH��BL�]�c�.��;ӟ�L]��2XQDȎ���r{��	��h9�{�$��τ��5]:�)�=!Y��!��n�����v���';��y@�JB��V?���/L�E?�F�O���yS!�D1t��."ň�M1c�d����l�.X|i�7XQ\��o�шE�TF�t=R�V�Ur03���ʋ��)D��6�K����ѭ�g�}�?�4M턻֎k�Ē��]g�-�KJK���4�zU3�6���Z�*��m�w�r�G�����C��l-o�4���10�=�ݻH�}�Pg!��h��&wۡ�ڦH�
�Ʃ�W�k}d����\-Iݱ���0g�a�&��?Y��Z���`�PD�n[�$�%I��ř��y�!������Ov�F�{ro�H���0h���s4l�w#�Ե�	y꣒[=�Nٞ�@����^CC�"u��ZO����!���з'�I�	�'�_���v�}�nv��sJ깞�)��o�Z��n:��Z�܄��`%��%���3<o+9\x��D��X5�=#(Q0�{+oV�v@c�z�9$�p`$��5�� T�?t��7���+��E=$�{���C��g-ƠCm�*��L��e́,(��OD�ɒ�7���gGu��3>��0��ѣ��� ��)�!,;X��K����� �X���
�f 3 ��ϝjM2kbi����𢲋�f��=ӐC}���"j���V��E)��5�K
��W��ڱ�(��S-�c0P���'�*բ��r���|=3D��� V�$@�%?��5��`�CRu��vf�D��id�z�uc6)@�#�3{���B";8}'�7�W�:�6�k^hU�.���3�7b�;RE /;�bH�n�קU�7�\� i��k��f��DqG�+}�qm��Ç��X\u|�,�ŹA��7St�;A�i�8�Џ�م�L��c!4[S��M�.Ւƃ�j�T���
\Їu��_��NQ�*�۹�yB�y`��y܃}��:�@��q�7#%���h=��K��p���Y>����%��MIESb62r�6�|��nR]l�|5k$ƢܦW����>��Uc�����&�Q�
�:h��YT��(:a�]Ms����̻���K2h��9(2w�PJ�n�5����<?��s`�}�ε*��o��4�#�y|��B�驎�F��=ءY�X�[%�}F�f���*�-����Sf��Qظ�Y��I��{4O7c3���>��������v���]���,��:|�m�����zň�m �lV�1F�iH�L뱜��������3����{��@ 3��$&��uHk�K�c{��׳Qb���YI�� ��u�ݣ|JxV\��t�"�!�&
ON�y�ʈ3p���o�9����/Z�s����I�T�3�cl-P�sd�����Z��Ї�9�z�V;c���B��w�e���|���7@]�b���%
��$����R����=�{wG0���{���Qġ��.��b�$Qݛ�#���H�c�n�n@5P�~	���BY�3t)�ыa|	/șe7C�G��$��z���i}�3�����;c�7�m.��pa�?�~�8ٱ��'$%��ڏ��g��9rW��}���z��"�0*�i:~�j�%����h��겗k��5��&|�
c<���r��:2�m����e���%>��ӜgӉ������X^���Kb
������8)a���b�%�~MTk�x��Xp��0���umХ��Pj>|�Z{���p�m~.�7�յ�<r����N:�%����E��z�wr������.��d؝2��\4w*1���>�	�}Q�@m@iK���oY���6������G�>�-���h	_�ʟ<oIj�Ϟ�St��D*!�짖5����h�님�_�0���g{�q��C����,�O<ŠQ ��$0QZ!@��Bg��*b|����Qe����[�ֽi�[��q� �!ej22C���*�^���p��N��Zъ�2��\�u�$��KZ�nZu��Kc`�E�T��z�%->�U�@ �tƥ9����G�<g��)F�`�� >E|l��ۈ<!��W��*��s:�&Qx��ƖZ��?�	�)a����8���|b��\"�=i���]��[��G0,i=m��:�b^�ݡ���|�VΪ�(Ρj���ư�y��Y8�6u5��,��e�������ǝL gn[A/y#�͸���3i���8�z�Ŵ����0��Q�b[�)���P;v�}YC�+��:F���zl�UZ�Es�D��
G4'�^n���@$u���ZQ���)�6����5��^�C܋����`bQ��}�8@�d�`��dc/O_YD�W_�{X��򎷗�f࿰d���Y�{��"��a[��D�m�12�f�y!��j�VW� Cz���:�;w *2\C��G��m�����Gz�,�d"f=(D�k��u�6���s&�4z� ��{ g@go������� ~n8��O�$5��qF��z{�����B2�%T1:b��W8!f|ח��BEM� .�#�(�҇�t��޶�5��Rs���og&f|�䓎���S�`D���ْ�!7�>%ma|j	���}��H���o�(ɒ��ܸ��~�F���nHk��,H����GLRH�_�V�K�iD��O2� �w�\k�>���[�vK��=�G�����������^�U�0���a.S�0�fv̑����m�����k%�S¶����F$O/��Rp��'a����xI)/�h��ާ܅B� �<���]kA3���,.�b���NHi��v���~��	-��ưK�7k8�̎�����iڪ�\�Y���{D΀i�����W$�ۗR)���s�y�	g��F�s�6ݝR�@�(���ܞP,.�q��p�=W��9����;X7�����j4�9D �F���SW�e�ap�\����lM�^����5a\m[d���=:���}�@��Ei�Y�ɏn� �T�����x�/ф����BͿ��_�$��~ȦV�pq:g��,>i�Ŷz�*��A/q��Qz��V "��ރ��|�Hࡉ��p@��V��z��p�0�� E$w�ݥ��:*Vh���+�~�S����G$��t�x�n��n��[�~�z�Y.�v���B�����a	�ϟ�|�]s�]�B.�����fxL�Hr��a$.\ �P��Z�
N幠��v�}n��І��C|9�}q�P�M�H��s�}KH6���ԗ�z��"��դ�
�ڑ[�߁(���⓾��z��V�֧2���^�q�X�-��`U94�W�[�x����\�*��k��V�4�'@øQ����h<��r:�9�f�Ç�h�������,z���$�-���M�_"^��-���mX����������Ւ�Bwض��a��F~"k�^7�5�7�lL�1����,?��۠U��a��7���;,�Z�����+f0������5��?���jT��SR�Iq9��-*��yb~��}��\��52ߊ��јa��Zq#�X�m�5}[>E��0�3��G�@�G
Ȯ$�y�Nt�_��_���Lmj�sSV,6�ޚp	�m��K�2P��* ��#|Z������:�\�1v�φw�z���0��c��|�(�_��Mcc�|��I���vk{9Y��/ "��@��	�N`xEƱ�^Ą�@�Gf,�9#K{!�o�W<Wb�U9�=Di�-��U�J ���^���~�*,Y�L���G�W�TZ�4��
:j�@�@��7ǝՏ����V��P�K)x��^�Rg1s��YD���R)�O8�;G�}�`�� 2��ư�]P/'"3Y���Fư��XIV��l��]�)7{�6�|�φn��Y4H'���K%��#��c��:��'��~l��&��0�Z�^�:ߝ�`oC�vU�*����a�����0���Lr�w	��p	L�F���,�y�H'�4��| 7C/�8$�l6����Gr��.�yVļ�C�E�~��4�CV>�x�lZE4�WnY�����j���g��4�b��U"�t�z��ʁ�����J�����;�Z��N�ֺY��~��e:��k{�0�B��q)�w<�o�U��Faku;�f]�Y�	�� o���s��]��^7C���j�04Ί���o�Lpe�>S��QJ�d�U��!�@�k���>ܕjU�nܫ\��fÍ�6�6r�z��w]�f�D�
(��՝ψ�MZ��)�uP'k�SdN�Y�O�Q��ѧh�3q;�O�� �;�]�}���q�|
`e��?���Tܤ�a+���{[.p�f��`��r���T5Wx����g��%�����W�Y��x�5��������0���:A5����dq9������������_w�Q!��}�O#�2Z�9C�5#!*���?F*�0cu���dޡl*c��I��h8�V����oS'f6��JU��p�F���r�'�EGZR�����y�#�u�A�3�Q�f�)\P�!���ŝ&J��5��ꆎ��EZ[
a&������d0��;g�U�\ߥ���}߽.G�k�Ԩ�B�~p;
�z�L��'�M׫~����&�a��*�K�̳�'6Ü�0��gtU-���0*�@�\Y~�X��5���
K�`�ߪ�4v�/�"���R�(Z�X�����~M��f��҇r�6j�^(��� ��Qr���6��v
���V�3!��zH3^�?�L����U,1vzY���eѠ͉�x3~�CT{'h&t�ko��-x��)��:@�	��Ӄ�q~���,E�Lz��X�8Hd��I~��]��G[�{��	� }�o���Vub��\����gD]c��Җ���ˀ��a��7��,;� x�W��\����辄�A�̷M���PWM$��@1k�ҁ�=�:���r��wE��"��Vp6���jɀ|�؀����R�l˪�u|�J����O:��ȿ�3sl{�����O���;�]�\��-�lPV���M���<&CMO|R����t/�.�U�&V�c�j#;s�U\��������p#JC��Q�3P����!��ߚ�#7U�ղ���>�O�������u!#</�����0��w�"��{��!�X�&��״�=�WM�`n�����%�*�1`��vF������!�R1B���E�J�+�(��ߢ+߼������9�������e�&4=��à���K%��s/�i���<y��Ηg������Z��IX����]S���5�BZ��2Z{
*3t������S$�~� ��k�+Ե�i͉V��J��.�hQ��[vG�
���uj�SiYarX�|�`4`�]^��A?�O*,�̺Zr�N����ܙa��r�	.��7�)�~�O%�+زx����|#�cGI��Em�q�G=��g9� C�nt'�s�!�L5���|�5�~d���Pt#G���eŲ ����Sr/�L��q��|�n�ޠ{څTR�F�鼸7��vK��`���m�i+�3>pQ�OQLp�s���[�ʋ>��i8�J��i����<�^�2Cb���2�Gql���ˆ�Lyx�UI���n�?���?��C��~�C��"��yRYu�L��d�V��ߗ�]�:��>M�iU�
Av'U!uVa�k�����W��oYק�Ƥ0(�=0�@*���!���v��Y��I�}��+�O����bC�5^���QjQ2�"�.��9ߛ��_R�XZ]uUDy='��l6����#t������p����.�
0��菊wԑ5}��|�K��K���k��Q�쩈D�ww��x6�n�}ǖ�7z�(�?!@>Хv���/1����U�h ʈܱ|O���p�9W�З�Ԙ��NLQ�����k��"�t����]���ZR�����Z��j�/�����������>u\�z����p�q��x�y��շ����/���b*�'7;�5�V���Fw�����>���Z�}+1�Yj(΍^�Lm�l��}Y�+r>o���=ӏ�q��$C��Y�T(�r�h�|�iE�e�^��tU�C�O�.��HȨv���%!e�r�T���&n0bﶣfb���B�>��d!}� EW�k�� "3.(c	g��R�AG�V�4��z��ݨc����+a���8�5��q����8�ʛ�U�����@���n/�R�FC�Ai�{�dePk��_���	����GT���Q@�2�����Ԓ`�yO���]�>�?�H�}���x���@t@�X�{7�Rq� y�+(-��샿BS�v#*K��*�%�G'̞�h�a¹�|��C�9Mb�]DY�r0��jN8] �`��|��E	
�	u���UU��tW4_dO�.w�Vd^�%sd�,���6�o�)�� lSmxT!������e�?� 6�c�vw޴c��i(`�V����˼���	ze���sQ��Z��:	GX4����xޏ�~]��-���;��U�Xh66��~ ��IFV쒡�1����hsP��{�1����hnA۸����81�rIK1���)�O����*������Ƒ<)���¡���`���ao?T���&#߬�����Q��[#�.�i�MLB���L��v+0"�6;��ë��P yJƪ\#�5]P����4�YW$S�I�=*e��d���Ƥ�?��5���!������7��/]�X`"k�\�b+���ԍ�S�Wt��Ea�I����Ԟy��ή:��ڭH�T�b�Z8x�L+�%�"&lZBO�0Kqb)�bIp��C�v���ե�@#�ҼOE�}��1�0	�s��Y�(�AK2��m�x��۽C	$����j`��gyl�]�=g0�L��D���g�����'�U����h��]$2Z�K�j��	�P(�6�C����4ʔ#P칔�JMY�*��Jr����/��|V:�+u�n������ߝ��VkG���@T|
YvC��G��&|���S U��{��e�n�����i�(�d���F<!aݮ�^��{6F��x�Na�g��Q��$�[�3���A�j�Q��w��ݽ�)J�'�7�I(�ggMi���I�蜳}�6�Yd���2u��5�0j㦠6�������X�b�X���k ep�&*�R�E.�DP���z����:�A�σ��l��^���<�.���շr+�f-�A�lq���w暳��|�3�q����
���7�1�h��#&��\�9��w@8u�]��j� ��؃�l�u���:�b�\��<l^5Y*=���K�䷞q6')
�:䪋�X3��$���Z,g18@�P���{�{`�WbS2{�A||d�(�^t��-Ud��z�o8V��uB���T���`�rX�k\�8Q�U��S���D\7��u ���2�#��e�����$���rP�+y�?q��Հ%�������{�5�o���}�s?K���Y�D�HIB���IR�_�2���k������ 8V�+)�U�q�5����x��v��f�[y{9yѳ/�v�t�:�G2j�����Sa���}��,U��:������1.^a����lh���8��9V!�I���r�cR�p�D��@ʅ��`e�>��-�q�  	�����ur�}��>��9��9��	YKSb)CS.3����0��@������P����t�*��Q�E�o?�V�8���zDG�%�X]7��R0��^ӟ��e֌b�.|��FPlEu6��Dg��>\(]�����N���&m���#(�tRG�6�肦3����-�������L�ܠ�y�}�������n3��k@�s��[r�{G��_l���Y{������|� �/�L��m��ܢ�~p$�W<O��f٠�߆��+4�jk4�R�� ���Ȫ�!�	���/��u��6�r��S��>Uq��ݗ��6
SO6�jO\�el<�==�2��e������^�xx��#9�#��V53�ʤ����u�<�`���8�������Az�����;^36%���Qc�&! �ȫ gwH�0B�}|"z+���W��O3	36rt��E�N�"T�](��b��˩c�t�yri��ذ�`a:�x�h�l1<�d��~>d�ؽP؞��e���m���ʩ5��b۸Ә�O2�B�숍d��@��8�a��l�r�wf+T����(��$�-F?)2^@pa�#�Z�mA"��g�X�W�"��$�ѽ�����8�-#����Qs谖|��E��� �;��	���C��_=F�y�Ϻ���䇀�]a4�ă�(�Xc�42���w�-n *�'ۻOO}2A#Qmx_��v�B@�e�>Hӛ���gɬ�&��o
�X��#Zz�L��_������HMo7�������n �)=���̅���x��X9"W.�xwȮ����I�Ij+�H�E�1}t0�0ƭ��G|e��E�X�]̀�Y^�� ��v��K�"��(!��\	^?J�%qGmy,5��P:��X�v��� k`4�;��;\��C���_�퍤�*>���$p�7[߂_��\��$���ʞ��	ž��E��j[X����C�;���E�i�u>,<�߮S�*(�"T[?�o��R��Ȭ�!���&��l���%��e�m{�M~�<s�4��	KR���9�n�YR�}��j7��K�,m@҃�Ӫ�DiKu"��M@n�?M_��V������z��'et����K{���&ʽ����Д���x>�SP�g%Q��T��
���B����+�W�0C��;���MP�{��_H ������L�H)�g2��y����y�剂M|����j%[(�NA��G �g�C�%��o$�]sN���*pi$l]��E!��rBu���z�S_���Im�P� �\ � "�u�Q��!�(�A���ԫ��M�X�G��ܽ��EB�}���F,�6=JF���p��âUJ��G�h�a}2��潗�H�Hkt%����j�$`<-�K"�Ą�U��G��B(p�W��h�b๖(�*����ᡪ.D���I���1Co��1�ɮ0���i�v�,��J�]n]��㞄ۚ�@�t��K�JkP�GFHi�e�3ʤ�9�z���p'YX��^ƔNiY�>���A_�Gn(��|�Z^Z����L����?�ڢb�m|��|n㈾�iE<���<�ޡ�u����� ���Y�O��~W����tq�Ԁ���.O�v^}e��-# h��o'��Jq�M�F9#�d��-7�g;A�*w(��c��:��ݨ@�*E*�)VE�Q�LI�[Pz��?)��xb{�r�vLT�DD+�~���}�j�v�|��M�zSYG&<�Nm�1w�D�����U�\$a�q<ӄ���I{�Km�_�-��/��g���m�1n��d)a[���dY�����Uq�ɾ8�EB�o[�������a+��@m"0��1?���'�]ՏI��,/~����l���)J��dwG����|��k��7P�^o�USW��ak�8��cL�'a
���X�FI2��_���G`�k!��4��Qhm����ǲtSB���[���ο�))�g5Ɲ��a!w/i�t��n���0u����[o����LWU�F�4Ր���� ��f��b/���1���ےp�b�*>�)���z~
�� �#���j4����uD`��²[���̤qqZ���^���V��Y��yf�d�:����WB�����%F,m��h%΀7$xm",T+���L���|Y|�~���md>q�Ӎ^�mu�۔5"���(>�Q��#}�Fd�߷�9l�"�
�Et�� �2{:W����Z8��y\S���p'>l�J��K��t��޾���ս��OEid��4H[�G����t�F6>?v�Dya��ِekCڔYs�Ԇd��M�X���q��}Q�X�˄�v2���YLĄz@?ޞ�y�P宨��H��3���B�,Pe���d����KiL{��
�ڕ~���X"�z������&K-�֖�? w����|�wǘ�ա))�l�~�M�4;��$.&�v7ʐ^�o��%$2 j����}��^��h�	��xӞ�RE{w�)�>�d-�wiѧ����_ܯ���6�f@Ys���aM}���@���y�0�0,�8��;	�v�s���!�[�s��:K���_���g3bO�Fx��\��u �n����ti����#&���%)�T�����:)�Ӧ���np"Q��:�Ϡ��}z�/aU��R��طmrE)�8n1�U��!;M:����廖&�܂Y���`Zl	���#Q4o�$b�B2������"U�Ҙ�oc�ib���S�Y5�EB�,ݔ������Z�2=@�/��j�E���ѤGXl�=��3�UJ���YD�O_����>�-�^Iqv�:ZyId0f2��A�0�<I�p؊.7����.��)�A�ڞ��<��v�T�$}�&ك8�_ ��.��m���5�qT���0� X��z��&�-�.���^�d��`&�㣻�?�A��u�:STɜ�Bݢg:���`���u[cs�����@<z�>#�����f��];��ԛ T��9\�|���%��z�'�+�S�=���S�2��T�,����vh��|UUU#�uk(�H]�ң㭗�7q:M���cE0�U�Ϯ�F��n�	T��%�Q2`$�hr��l���q�3Y�;~N�b����<��\��غb]�s�^�YCW����ڻ����;!7̻�n2.���~�ߪ��llH&߷]OE�,����][βy���ˈ�[���+�XF���wc+r��Z[QzW�-(��! ���m��S�e׬�P�\U�'ޯc�=����H��XW���(k�����\|�(�/��J�(h����ؕ.IN�@!�V�Τ[_������%N������ﮐ0B#d2�j��,;E�qjsb��lǺ��dѴR���n2��.麌
u"����m�<�l�T?|����W�zVB�O��¿��v>�)���/xz��Zp�����jb�w+!z|��A�@�H�]?�3n�+%���u�q'8U�n������o��Dk�7B�M@�m�����\��[O��9i0 ��3m�>Q�q6o��%T����@��u�+L��S@�b�!#�y�]��ҒQȄ�������_a�I�f-Z�4�5� w'��k��-���n��ǯ�f�;�S s~^I��ne���+�	���)	Ĭ�q����W;뱝���өP�(���E�4١�͂<@2���8>eB��`K�mrj��$*�!���l����������N�Eݎ���^���wPy��OL?�������GB�0;�^L��7F��c��ZE����Ԩ����'��v��iᅩ ��&�>�.��@L��Lg��X=�P��oۜ��&x�v��w3��~؍�㤫i�eݰ܊y���D�k���&$
2�?�dLƹ|��5��1��=��VYs�[s̮���[��$��B�Q����������dh����n�Y\�`,"�3y`�����d��mH
v���!t=\,�s����_N�p$	{郑C�wo���J:�Q7���b��6���FGP�A5Jaz"Ϣ��@%���D��zh�q�YL��E>�G�� b L"҃��iH� 9���U�7��,J�]�|bW��H��I���P�T3�ᄠ�םб�<�/4�?���~��z����El��Ď�F5��Y��06���
���/��@��P�gWZ��pqϣ��w��1�X/�3E�'�d���򵄺!C��V:���uȳ� �M�pUT���c�5l��^T~V\�)&�^�#�l��ϼ�d��5�~��˯��_f$���8�D�PE��$Hў�pT���LQx�~3ۯj��B��s�v���t$[�X�R �@�g��HM�������n�ǰ����Y�޳
�m}<� %*	��)Sm@f�3yL-�i}���y�UR��>���,����Xx�q-�quY���g
��0�VϖȲZ(��~�Z5Bb�x5��Ё�d�,cT�*L�~mB�xƊ���QD{9��NJGt�\�5ϻI/��l�̤�)�l.mO���<uyK��~b^Y]ZqL$�у8e�F7V�9�3�v��t�&�c��d9�h��e�2a�d�x�J���/�e�ݵԕ�#�Oe��|qŹ�z����8r؃ۥ'D��	���_2K��,T"Q��5"\���
5�r�۶�17~ͪ+���0j���X�V�$��!��̑s�����5�.nB͔M1�N�`[}`����2��R����)T�]\[�T������n(�2gѺ��G�GՔ�˦+�(R.�p��-�?ʋ ������6��lZ=����{+��8C�
����WĖh�ɻ~�E�Q쥸`y�+�J��&��;���������wj[v��Wt���J��Ba�c�jf\�٣*��2�V^j�;�M:��
.�����nϔ�9��F|עc�u��Ы�ޞ� ��[>3�=� [�?�r�Kez����{�<\��d^=�BΖ��,SϿorz/�md�%Zv�P[=��P�F��-�{�SS�uB'�
3܇��v�Wz}��� �� ����-խ�.�!�q����. ��k���3%�L�CX��Z#�1�������43�� �9����4���kba�:5c��5��=��;]5x?���s�����՝G���F_�L/H�A� d�&˜�� �n�7�F�����;��;s��e�&�(�jQk���t��
�fR�^:o��t��w��Ii,M���1����M����Z��lZ"��m� $�N[ ��!v�-x��m�(���|)�,[N��Nh�b�%�Z�)�j��b�J�9h�T���r��\�T�jmQ-Ǣ6&�Ev�/��{�.�d�Vʾ�d�t�޳�q�[����s�=�"J�d�@����R�.�}:"�k�(��M�K=J�q�ː��R���f�WA����{��=�����?�x���1T'�Jp1�"p���i�#�[(^XG&�o��2c���t�ʴ����nc�Y��˄t$1i�XV�ۓ��3�,G�[�*��)��o[ �b{Oj�S����I)J��5��d�T:.�Q����*��M4';0bM�y��TՒ���;sj�f���z?DyR�QD'gȞ�Pq����?�K9�Z ������ײyKu��?I�t)����/H|�R���VĴo(՗T���/nb'�ٜ|�x,&Ձ��[SW�^����{�X>I�� �n�O 9E�.�j=/�Q���Ǔ�	4}G,�}���|����.�aQP�@|N/HCc^�[4�Bc(p
�]E�C���G��[�ۖS��wAqF��QǷ��YBj]��,�-o��{*(vGm����$ Y�-�3�gв�u#�f�	=�r~]���B�c�_9�� �4��]9���d��k;#����ԄNe"q�&M��/������n&�*�6�����=��L�;U"��x���̴4�M�}���z��C�/6��&�YDY��x���pq�BP�rK9MJ�Ѓ��?�ꍬ���`�.m٩q%�aS"bNuHx¢��]J�j�}���Y�b$���u
Z�\��_��r3���t���!ISU���a�(���)u���4�8:�'��%�]1��vL��5b/M�Sۃ��3^�\��G���Չ�;a��`�o�	��o�޲�����K��i��!��W������ɝe/$�).\�~]|�.��o��T�CJJ /��'��y��_�m��Ġ���Q�������$����.�
�
�yHD��\�Rs� ;\���8Cj$�c�[QH T䤨"fTp]�}q0����+��6#�F{A����J9�$��C%��3ۍ(��Ί�:@���a-(�S"ۓhWg�kta�6�#=�8��(���$��V�/4����*�xa#rVΖ�^��܈�2�.��mn��}��.��o�`jFh�,�g}ʜ'��h҈>�;}ێ@����+��\��5ϧ�~|�Y��J���r
�բ"�}e���Hp�1��8��я���(F��L��e��z�j_����/|���#D@�n���$RJr���ؑ剏P�3*�(��V�76>�Et��6� ��;D��)d�^9}P���rQЛL�p����JF�����~��F��_�u5j"���@�"��e!�VN8�/�A�ئ�]�X�F�`���_��X���x�^#w��ۋסL-}?�@�y7�:h*�u��X������t|;]4m�Ml谦����@A1/A���u`��H(vVGZ���bsvR�$��3ʨ19�&	�fW�no��q$@
>#N�#��q�6��Pš1���E�jQ�Df������T��a���bSd�����P�N:'�ѻ�~o^�ph	��u���'\#���u�&O�l����Q�5���|��Q��7\,W>T�!�0?f��.	�m?�
�o�P�D|�ײ�XĂ��q�l�vN83�5T��B@O���)��_1�$����I�*NsYoi�H� ����+^'"1�&�o�J��%�(�֏�]m5�B5���b�K���l�H�����!���r:�ר^��l�LF%G��c�;��b��bߞ�A��B��8��r�C�I~��H�x�
���ܤpt��t)�m�뛙�x그&���ѧ�jV⁏g����� ��飫�V��"t�P��h]�1�c�G/��[a��6���a����BŦ�w�@��
$5b��y`2��� ��i�O\M��˥n�^���Q���~���!
4s��f>�%p��16�Q:ý�9R�$��XiOėID=����"M���1�����A2�o�Cca/������*Ϧ��ۙ���Q�E���-�D�qhc0Mt9��\�A͉P�!�lwI�?���o��o5|��l�I�N�,�0�?5]�����2qt�����i�zz��R��;��Y5ZIyދ�ݦ�0�����c7Aש˨	u��j9��ȶL�X���d�U-��ga��˺�M�~��
Wi������bm:I[�(�� �0�C�c�j ���vG�m��i�/�BQMc��h�*S��"=��������R��ѝa�n<�����0L9�w�~{�x+��"f��Xu�� �!��əх��׏�3��@�)0����<�u��X#n����4ob�J9�3П���V?�4���J)�(�&?����hxT]�e9�ڜ|�ӻK����t�";��	�h�ڷrs��!��=��<�g�7���F�,�E=�-q�����C88�~�X���+��C�BchN�թ��H�KH����a��s,��6�9�If"��k�s>���?��t����D���>��kb�1T�	_o#�@M���|y���Xi�l�����'����j���i�O�6b�2 ���'w2�-4�f^q�k�� \t����Ϝl�����,�N��� g������=S�	M�
�����,��>ۓ�������ʣ�M�Մ����w���|�dncL�^^�nB�� 	��`!�J򣢄]��څIw��n�֜ۆ�6*g��;կS3r��G�ǿr�]�ÍV��{}��#A@~6�f࿞;o��_��˵߼�c�[r�V���Q��9nG��\�[������O�f��t5��m�L��r�s��<����~��M؃���b�9T~c���5���w��o%%��4��I�l�y�	���!|�{'�~�=>Z�P�{�����M��ʪzN�*]A�f������,?����2K_����ώc�ξg���֥!Ș2I��y��Q�%���XR{��
 �����j��Q����Y��1Q.���'=�F�)؁K�=��L
1C������8�� ��z�VJ{���t��f]�-�V}���25�����I�C�8�}-��(�V5�:�� ����@&��`)�G>7�`i>��,š	M��X�%�1�:s�U�k��{
�:�λ�
3!u��^�D�Zv�.���p��^yzF�+GZq�p隯SJu�v6�����gI'�����P��E���������B{JE�z�ۗ|;y-s�n�2��'����=��zAM�0A�����/��FV������O,l��;�JϦ�1u F�x����s��\�
HC���I�N�*8Xt����o1��G���fF�Og�4� �-��Mo�-�o2C��U
H���=G����XE�{�6>�a ��K?�������v'��
UM�n@~ޔ=t6��]:��0䴉,��q��\V��&A��������=���3mF.�`; x�4�9Gy�l#��hi�G�J�,[��.t2�6�kȱj{ٻ(��/}qb���Z���X�9�m����X�����o����� MI���}�Q�iT�=��N�r�.m���!���0h��Oo��d�*�DR܌���]�5&p�^C1S���Dc�q�Җ�ӒÇg/����*���X�}������(K�%|����g+���-DVSm��'�	؇-����WP�W1f�T��<!������=�;ޝ�)�X�|��*�V=O��;��wMg(��z��$~T�ǃK��&щ"�pºj��4A6Tn�]>���}���s`�/�"��8�f��u	SD�X�Yw�άQ2݃ CV
�(}�)0τG7Ut�k���Tx��U�C�T�8���؟ 7��B���,�'/4��+*)�P |��U�mҘy�:�=��$�5��(W��l�앎�D{�g��rښ�$��6ު#���h�����R�8	���T#�(]�O[��W�a#; ��ϩ��c�ڞ�aXwܭA���[�o�BΠ[�J��JD�}e�\�	SiV7ʱ��I�F��H��(��n�x*س[L��{	�PpL�<��tkg�5���f�d� �z1w2���m��Y�bj�D�~�K�r
�IT���n�J�! ���ׄ�L9:�w��X������%�Rd�I&)��ވ���B��w��.`qWk ��C4�K��1�Y���$n�V�y�7}ε�] g��^�z��L@�\���LW�<i�{7��y���bc![�N���?Շ�Fu&���K��?P��s.���c4�`�@�P�2��­��E>ؼa~4ܳ��<MQ9H��ơ'�qF
$��2(�K/����ޗ��t��G%�l�t>�qEn��T��ũ�=�=��\<'[��؊��i�$���[:�rob���A�� Ub�bS�d�5۲����H�f�=�M{hc>׀��|+
���G�L��z�L��h$F�(� |�Wo�t�wlU�fͲKH1��Q�Z�w%6g/3�(7�C���y,�N�)�;{QT,S���JV��82��[+R4�^�w����?*�"���'ޠ�n�\�:JL�fe����vp�^D#İ�E�]����l���sG���,��p8YK����<�:C�,)����a|sV!��/ǁ�1Y�X?Pd�,i��hz��sQv����>�� �_)P��$S��lo��1m�h(d<�Y�it��<u��aM�e�3�/i�ȗ����/���#ƴu[�beY��}��~y96{OM.�����0��kgLcپ�~0��?�ʱ&�r�L4�:k��@��ÿ�������S|y�ȡ���L�Og
P���b�6��-=3���0x�a@��ז��*�����t-��]� ����᝿i�G�ٴ�Wϯ�����k��r6�/��O���<3���XM��	9�&l�Ɣ�M{Ў�(l^�鑚� �Ib��MP�;eW�Ϧ� 3�ZGHg��.��M4��C�n4_��^�A�5��d"�Ȁ�<R���aIn�R��:��Z樂ӧ��<���;�^�{��mn��$[��=E�<h�t���{d7!m�W��������_~�|$qG�^B�R�� IB������grOF��i�abi�.SC�7ץ�NTj�S�r���!Y������,�12�Vi�S�ק%�M&��ZA0��C��n-=�,�G��N��udk�dN�񻚝�o6�-љ��K/��.1�--�����$HIӆ�@7���t��_Q_���	=�~��YO�<�.��Vc�E�G�nV�^�AW��u��8,��䆺to��I��y�J�9s>pS��oUۧ��b��=��zw�Ƅ2��������1�P9,e����@~�s/G��NDP�G�.��:n���zT�ja��ES����͌�0���|�쏴-���U�Un�ϩs�*�b��:@T�nR��a6�9�8rX��J�>�����#�h)��׬�e��8���&x�_@OS�m�F�|3X�TD�#uI'�ms�Vh�B�^/)��"�֓D��97J��C�lB���+c��KnCl%�,��ʓ��ֳ��Wȿ�5~�vb��WB�Þ��S���nE�e�y���y��.Q��7`�&SV�AN�1����6���a���4	'�-��5��E9���f���Y��X�yݏƂn��q�NM�I�KȆ�y)���L1��3�"��t5Vz�"��,�k��ߟZ|�)��*��چ����<�1x�� ��TKǇ��Ȥ�ZӜb'���Ln�<�Z�l�BZ"a��.1��V�[b7༙��X����>ܹW8&6���W0�m-6G'�)[�wb*Аc�]�t������z.�2�`QvQ�8�.=�t	hDk������	I�T��"C�o䌍0�,��6��eO�4X���7��ۧn�8����s�l���H
���*,`�ݵTQA��ޙ�B%�ǟF�4:ᜊbq�i��ĵ|�=��&R��Q�mBWǒ�@�S��&!����B�����.TF��&�<��v���e��s@��G#Z)�c���:���$�L¸�T� ���@����b�������E kI�l*l�+T�0���xg�J*� ����N�z����jsj�a��n��w�R��&(�['%p��yO 2*Z�`M��P��,�U��=�A��<��7_]��Mk���xj8��p����[�����aJ -y��O%�v��z-��19���UbG�<���o��<YN/j�wz��\��[�&Pe�,f�w��N/ �k8_���3����5�1��4|��Z��8vgl���D]��r����K4JK�KC!%��;(7��bQS �y��[jj�UEz�1C��.�*���]���=��/.��Ǒdy"Rb��E1�!%0��Ͽ���[rj�1�样�@�I! ;.?��:�7�4���yz"�D�s�ϱ�0h��@x��>~{��oP�V��M�J��M}{���S��cJ�{s��1/���c@k�ȇ�=v<+�k��X~��1��$��W�����C���6�L�^�z���
�W�����`l��%����'�r�t���8i̫��I36��h�XB,,�4Ӑm���p���yJ��*C���]�gr��T�K*
��c�֟��a�b���xߓ�����/�$D�6.!~��َ=.VȣkM��d�P}�kJ�%mg�l���
w�-�O|�ծ0P��̹1^n 0ĥ�J0�^��X��.�r��k��]s֧UH��uhU�)e���~���r����Ljy���y�����	�-r��� ��aF4��$��(�(r���Oe5H�v2,��D�2���;�g�#�J3��D�����ei�y�LMB&����ڮ�%�����񰙆b^\�A���]sZ屄.�	u�0mR<��q`�%�O$#��.�6��J���{TU��+9:[`t$QNˮ�Hn�����.x �K6��O��B�*W�$�* ��	\��_R���Α�B�H,/:$lU��7z
��Ȏ
�4}�O�f�}�(=C�;�����
ID��b��]�ƹ��1��<(`���z��*����p�2M:�6��O1k��fi��Z��W����*@������;�<T^��te�60fǒ�Y+:fBǥ;x�o�\��i�-\����1��`���)��rqP.� Ss_0��S�2<�ᳮ�+1�94t�!}%�,� �3$Hҙ��mמ�	
���^PȺ�7���d��0��������mPJ��z��S�ϕq��N�2�3=/��
�y��j�H�3��:�K3{(���[4�S*xK���ʈkC=o�vf�5�4ѹ��$Ƶ�>.��5T�/�ܣ�_�걕T��0Jׁ�e��ȱ�P| ��i����AnBɪf�+cwk����m�"���Ρfo�G��I�����˘��t�ŏ�z2��/��@��V�'���Tp]a��+��|�P��7.u��P�%����F}�t6�Pʧ����4����T$��J���^ݐS�X ������)e��Ô�^�=��ז<���I����{L�UKn�����P)�ޘ�x�n���jO�+/��T�Q��:ǘ+�����W�6v��DrC�4�;�k�sv�Z"����\.��)Byb�a
����ݐ�đk�IX����J��6N��b2��I	��ƽߛ�����=�6M*��G���L� sO�%�f�b�ڌO|�:Tb��n�HAb������<�h��&��\��5�ْ���ԉ�h����I�f�nh(��F������O?l��d��x_.��)��Z���y7s��B����k�X�(V��Z��L�ˆ���\���f��˷����+h��M��>��t8���,�� ZOwdx�M�+�p��G����4}��2�b���l�L�����̐�J11Љ��������3'4��VN���{hE�t�	���m��f<��J���Uoj��gw-[�T���L��A����������6�uLT
R�SS|�D5�w��q�'���� ����p��v��-y��L��xӰ��m�	$Y,]�HT��\�/���-N�5��� ۉ'�۬iw����T��RΛ0)�����)
����<���3����a):���2�v���)A i�Om6]�Y�GV���{q��K��/y��o�]޳P�!4P�2w�?��9G��^ߛ�M�[F�����M%A!K���En��.�*�k�r������$�Ԇ�,%]������a{�hD.������&�]I��l�O�Z,�:`S�u��|QL.7T�d���ɷ���d.��܀�)���O>���m�#�j�AO{{i�����ʿ�vի�=�0����ƹ��8�^ܗisAK���O �y�t���MI�>:
�j'�o��aCĉ����.Hc�<l&�W�Ơyzt�y�X����ۣ7'M�}�탟�n�3�Lq�9� q�|�aM�&�+j��k#A�b�Z˴m�T��!�=n�Pp��Z���Xw�x��'@Uk������h\D&��ʻ�Q��^\F	Ӣ������Kh�5�&��:U=� ���u>�9Dfk���k:>O*[4��)�˛��<Մ8�� ��,�G/¼�FrDnf6�!��ҕ�L�"��!r�4���F�U6��Ƿ��	�Q��Ȇ�� �+밎c�&�[�'��A�_0V�^r����ng[C)��"�Knv!���Hƶ�U��2:}���7ժ�s��@Z-@����#�)$�N�C�v�Ń��B͜X#.�5{C�|Tɀ@zJ	���Rd��0��A5�
w���]c.*��}����7�I�m��`ÖD���4�g8z��l;���Ͳ%"8�"q� :\.�<�;U�7[Oa��݌D��9vy���S�B����<]W)��x����O���5��.��E�ƣ�I��p�ࠌ�4I�R�wB��b�0���i��<�;W�v8�0{*�Fke��3%���R�Hq�xoڝ Ɋ�lb>����?q�E>̲�~:!Y�8���4�͝j�1�G��+��5`�9b<BCȘN[F,�d�iO+VO���K���&��&ȩ�22�UJ����o1|�� ����1Q;J�_1iS牦�~e@��il����W����&w���$鱪��&uC�z��S��a��R�kxKm�o��($�O�Udi+礦6C�*t1*��v��t#�żi�9X��-ί���0z��x*�ų�����yX���h��D�!9��@��봮�}^��gɘ��_,�4�� \�(R���o�
�/�%S�*m�s��m"!�C�/��5�?i�ˢ�{�e�<6X����H-������g+A����C�5�X��K��]�]�Wjb5
�7���ON4������z��F��A_%`?�,��K3�	߳��
�ݺ'�������J�����v��n�5�C��SZ�&����2 �m�0���P3�Y\��a�,@1f��!�a��Ξ���97U�Q=���Es���ۈ������r6��X;\�I����E"�`3��ܰ��W'��������agȋ'>�S1��.}d���"�N�C�?1c'4��E�,��n��o>{!$�����Ъ���-o-�}��lԮ�qhR������~QY:��Y�O�;H�A{:+x����"}+�x�x�#_&z��'����#)�W���e~]�W��{�8��a�Z�It��T�w�/�B%ږ<'����'�`����"O�P��Ԟ�ޓL@	 a2F�j�>`�#��y%���#nN3�������n�Uz�D.	!�i��ԯh�ڋ�']̒
"�t�o&����.�͵��:�r� ��Z��Z��55w(��x�%��Q|�1F� ��}Tf�)[(+v� %!n��\bգ�o��S��)�^�M��5E��.E^YH���L���
0���������Zi
��F���u��Qi:� ���̒���6�9��ދ�I� 5!�G�l��@�hyH�M����>q��O@n.?����<i�!r�~0:5O����y�����񍐃i�W�לHW�b��J%����/|�V���f���.���l�L��ӜEbbYe���A/1#x�lJ��;��p��n<K��R�^Ž{���6��N���o�h�����0��%���������T�2��qiR��e܆Ɋ����bP*�:Ź K��.��!z�Ok�9l���W���V����G�2Z�>�'�,M�T�w�Ģc�=�;���d��7�j�z���
����c2�*�{�T+�A��	!%#�t�W ����c2����#ܵ�ZNłdg9#faT3z��X�J�z�����en���8 �Z-��'�㨿��G���+�b�d�~�}�i֞V(�v=e!�@����yѳ 8m��N��	!�(�' ��l8���`��`���T�]x��cC���t��;�!�~D��e��0]a.Lg�}�١��Teh['1��b�G�7�d�����a�!g�9ӣO5���������D��06p݁��8d��o���:[��X�6Z�v�D(L\������zpw��)�Y�M����d��������
���/�-�>� �t$Q8'>D���, �m�>��*�����ᚦ��^?`掃w%Z�n�5�5��eݴ�� �k3��z,R�1��4x�Q�P�qO�m�� g�2��x�j�կֽ���1���%R#�i?�^���F�{z���XYԘ��{B�3j���3�����~�B���ˎM6 �d�PK7�y)�
�W�~?)�,6��R/dS퍞g\~k��O���b��C��I�żI�e2�V͝c���&	|��������K�8v=�w��vrP�q���3nɩ˄}$�O�^SO���#����XZ�%>J6�p�ײַ,@�^�n�JQ.��n0j@�#gϚ+����_��E��!Q�5T�zZ�I<�P�'���+�� 8o,o���=̿�\K�m��k�$]B8�к�S����/���~Y����4BBs�U��ކ�1\��`j��"���a���8�q�ۮcOb.�נ���W��6GDAo��;o��O0��3s�<�hd�Fy��P����-��9�'r����Eb&>�u��F?V4:��,|�Qu[B��N�;^j�sK�mNP�5CO��3�uc��J�Oc�1����^%�i����^�FLq����V��l�]��s-(�%�T��gùV�v���e%8��[>x��)]B�5b��5��M?�5��T���r'����@2����Bq�h�G`�7�/az"B��e���m��8�l��1� �/�o))���,q��ԟpK@��X2���f�rŠ$G*6�����)_�񓁭��岿V3K�UҾ�V��٤���D�Z��y�K�"�Ac]S����D��m�c�g�c�G��WRVF�����y����5��k�ř�PX����RpA#�dg='>����q'ݛ�?�O���Iwj/�Ǽ��Cה�/�%q���&ʱ�d%�B�����6T���t,ϥD�y�p<��{��`yѤJ��Ǟ]޶�7�۷�����%:�i��7Ӛ���i�q;�p�g�'�\=��xB��_��<]����9���T#��a��0JOxǨ�8��)a��[��I�F:X��=��j.>d��Y�=��)�@W�H��\�J�1.!(�z^�����j��̧x���`)@
�����0skr\��#��<g�gA9<��|!�+�_��d�sWK��Y|s}�y��d5�o�tz���5�24oj9���i��5r���U���X�#hgJ�H� V�@�4S�4k�3xW�q]�V*4�K���<�Y���5ן��!&GW��b����6\���\zLB��ZR�f5Z\Kma'}�Fr�R����T����m�u[�٤��5}�嚰s�LB���,vt c�ì�����~��e'n���}͜h���Lk-q^�r)k�3��E��s�
O�j
�l�<�=J���5��ee~׿��/ث�m�T!�7��s,Z�4��R�I9:Ĉg���{{�|�?��6Ә���>���r�",vI�6�� ~TX��������a
��M�La�%�
��g� P)Ku}��b��	Ց�P�tX+�o%%*1��~�1�~�o��ml��)P��S�X���-�3�I��1��8h����Q��O���ۑ�-������z���_�d�AK��P�չ�(Z'��JTM��w�!�?3*������8!����M<#I�g�� ���\�+���Ce��q��I[�n��W���ά'W�W'z��G�b9�X�٥�k��Q�1�W�S6Umf,,���=�4L��S��n4��T�S[�R���i;Y�����l57�K�$u�(���<��%�����x�Qɴ���C����?>՜N��nre��� M493�kp �ѹ�T����y���!ӈ����q�X�� �]�f!P�_I�z�d��x^8��jĴ��r�I~	��(��P����T�Tr��Ă]l)�N'�F����m�y���O �0��@���A^��C��P���e�����+�vY�%�]�϶��[�T�pބa�ΠU�Sy�b��]7@x��t������-���)����J�	E�r�H�{�D���Ҕr ք5�?�nAے��g�Y�iD?|���%P� ��Ds���3S,\dp�������8k��.a�Kss���a�3Sh��>�6AJI��֒lGb'E�a�"�	������x��O���[j��9^�����|������:�@��$�<h�(%�6��V%���J���k��>���-�UxwF$xb�("�9�ѯ%u�����Q�Y2���(h�)@�� ��;:���:�M@��"q�χ�!��FK=]���R�B�5yk��~y�>��5��w`�e8_�L��uXKߋW����v��\�M&�lZ�\�v�f*����'lq�:/�t'N�Ƀ�3w/_xY�!K*���c���]�]3�z}qRy3m����5�0<�f�L�&���nV�@����V4M�ի�/IL�p`�KT�)�F`N�'������}��+����'��6<���=_ԟv�IkxA����/Wjpeb�5�߆
���GGS��O��9�A���_�(��Q �dgv�*�2<��*�[n�P�R�"|�������d�Y;�����7_$X�'��-#�$dF��)�����g8Ѵ�8į�����#t��B?}Gz4l?�!:hIݓXE��:"�X�����ČJt��V��o�K��, ��~s�z�sz���lB���?j����!�;˧���9��V�n6!�$/7�����!V.&��D�2Y��@�iXV<`��Z�_$��
��4�������$"���RSS�'�d�֡(���] ^�,������y�d�4�ݦ�;Xǹ�| 0�A��'Ul��WSя���	o���鿣���O\����G:]�N0�K"]��he	�0w���>��}v]mư&�� �͕���+#�3#hb߻��5c�/32�"�l�<���ވ�8"���lx�R�ϻּx�0P�8�i� ��m��&^���o�|6���[���ѕ���o��������hq�F(iz#�����K�tU��,cd�c
	���!VAd;(u=��ͥDJ�0���"��"����G����GӬ$s��֊�?5��TO�q������ds�^���[��dṄ�6���%�-d��b�>��촱��#�����#�I=
��ih��_>���R5�q:-�j����`�Pm�sZx�X�v��{xOA�Sv�2���&���5��]z�./-v�:���Ɗ`+�jѪga�)>����ݕӂ{��[�蜐�v� ���3��g$���AW�����q{`ݽ{��CD��1��g"�!"U�DQki3&t��$�[l��Op9�qn{5[i/W�\�W�i&�7��p��6���`A��i5�޳[�X�,�K6����҄b�~�Ux�S�G�D;'N�Mк#�v
ю�y6��3�l'�ֹ��Ļ��ӂ��#�O9�Ȫ�b�RNG�8�eU3��5oLԎ���Xs��i���"��K��w��=�M���[�PV���[�����ڸ���-e�~//��e�إ�g�g�����6ZJl�q����"������vr��v7=Hn|RG|S�P��j{�XfR�����2�����t���Q������uPk�f�(*D��v��RϷ��L~����Y߁��Tɩ�4Y��Fh���jC���L�y}�2.���tJ`Ƴ���D�R<$�U�̶)�=�;�3��ȧ,}Sw�v�hA�*�F�K�k�F +/-�ظ(�)��V�ivx��@����љD�;�4��?�.��>2���hJ��9�]<M.c6��Q8��:X�ڀ>LU�-^J��c�D�t̃V<�u��+ �W=���)��tyb>�s�[�	{2�|�|��o���˼��1_��|�J�s(�SAq�nؼٟH�9�&�EP��#��\)�����j��#�k���^�"���|���E����t�3ܑ��Κ":aǏQ�������/��;����,h_� �p0��[9cEI֨�^	J#�w8��Ր��;r��i{��#8jgL��۞�nZ.�L�/�vQ\�y���Qb�y��mX���aȢ,����"���ɼ��|�ٔ�l�G0�f�A�/����sL@�Kq��[A�B`Y&����fW�9�/o�,#K�
�9u�`��R���?��\� n���N�I��=<��G@�B����U"��X��B�No����T�c���;(X�պ�d`�3t�eʮK���HmS�?=Ȱcպ��q���Њ��ӵR;����mb�cɽ��a�MJ��F�l�Qi 5��#���mlx�<9qҎ�a�%{H$8@1�쿶S�+;���3#����P��4�(��{����H��/�Z��	�?���{���J�U1�sbc	���N_�ݏ�S����~������?&�RScxHƖ�y3y�?��r���)�����M1�w�݄��cNW�)��o��]�:m@T㒀��S���VO�
A_י<��'�Y�86+�����z�*��?�e���9doR�b���}g"I������(B,ȢOXl$t����@�� K�&�;��&���z=sf}dd�%��?ȢLq����P<q]�V�D�� #Fja�yZK���hJ��Ֆ��6�h�ڗQ����!A3����!M�-{@���y8 Y������kO~`�Jy��@���5-����b~��!UFNQj����W�cx8�$~O�>�����ӹ;�-��I/=v"��h_���*��ð���(��]"m�z�Lě�J��*۾�@���޻�J��^��B�G��s�)�l�e��R
�b��J����ݯbE��Q����'DBL��[c�b���:�4�V���Uc��>Rъ�o�HIi'���S�`��+`�*��PRF�4�������eu�t��x�X^��L3A'r,����F��#�Z�I&��V�N8(&gM�
�ίXQ �	���8�F �����#�x~ ЩP���q2��.�sS�Z=�7mp�WYf��� 糱�쁅{��4��WAs��Q�E,H�h���� $��7���Y%/�c��&�7�}�/X��w�g�L>tg��~���������Z��ٌ�����1��� ���ڳ	��Mˤl*U���l}nn�x�W��5ږS�D�:!V7���ɪΦ��j�Z�
�n�=^ʳq�I��O�%Hw�L�L�ȁ��%e�ݟ�Ui�7L�>қa=b���%!N��;k׆QG`�%D��!���K���4���mx�q)�>޲�z�x�xU\��{��[͘���'+���!ͰX�|�۠0wٱ��iB0�y�@�����$��B�;�`�(�p᫊gN ����C`��9���w��d4�[��i�\D�_=�mF9�U���0/��w�r�=b�E�WMV���K�t���D�}.��H�}�d�̆.��W��A�ʤ\4���T�_J l`r���Zi"��u�A��Y<AE���F����d͛�3�͂_p�hnT�y"Kw,�T�/�I�cqk,��J���ą�����im;)t��%@�F�4�/�x� Vi��Ɇ)�x�� w�n\�S�� -)a~�h�o�A̶V�ż�}�i=�Gw��Â.��9a�U�0�{�������7y]XbZ�`��	�~��4��B�ksVX���X�p�w�%��R��yc��ڎ���Q�NҋgA����@�ۺI<�ԏ�&x��{92�5H��!�jMZQ����[�R�i��r8�@ٴ�����xS+���Ag�g�&	��s<���w����Ȁ��^y�@,�|m=������P�����؆��f�`|�qE9(��`�"d�`C@����8�n���|HՀ�NTn[2@��/�Q͕ɸ������x�l׀�׆��CˆC�t;߆�@n�����?gb�ȏH�s��G�6ߤ[H���[آ=Mՙt:�<U���諺�� ��j��b	����
�~�*�����|-|s�;}��<KQ0�;~ϗ`�;����=�X�v��_,W� j#��gQȵv)�4x�"q5DiD�C�3�����%L	���&��Y������/�
������Z+�jUa��H7�@��� �iCD����%``���r�&��Ŭ��ך�#cdP{{��4�OH��r�b����u{ƚ��jt�:ʑ!*�y)����h_�n�^�cHY��\�\FElJCL�S7�禡/�s��8�Z����N2�2��ɍ�I�",�1�n�-_moֵ,DTtr����k!H^hҌq���G#z�~#�?CK�w���׭
&W�L9�v.�oiȚ6��[��TK�S9)Jjs�\g�\�G�3���Y��`�#�:��*)1f�(����G���:t,��j�.T4�Y��9#l�o���6
�R��@	�XFc��o���4�0�$)���[+���r���T=�g�[|��Ӄc��R�6ND|G�^2,f��F��$�%�i5������^*I�����STУD;w�溟4��R�'@6��ugQp<�f) =U�4u�s'F�>`�a�E�2PبA�~��'6����؋�`R�?;f�g��W8$��?��X�`�%p�����5|����ڭ�%�^(�:K�+'ʛƅ%�����G�ws�'PӛG;|�x�>�3�*M7���w����_�8���B{���ɞ1;��5uV�c�۽��k�{{���+8���%kT���Z��hz�lO$(��z������Ή1C�B�0�"���p`Nx~ ��Q$1e��Q���k���'�!7�|@S���F��n��������B�����vU�}�����:x$@�yT����w���A[nւ�kS[��%WR[��`���k��\��e�68f�߉O8eLDM�~l��v2U�, �Q[]��7-�jYcf�?��_Y���KD��/��<�ަ篁�#:�pvl��`/@��k��1 {?:Bo>6$E��������U<V6^����I���p���6�;�����gn���`�g��u,,�?�%B�Ҳ\`�7?C+�S_�����f��:�SǬ����V�ؑy+�%rt���H��h�+�!bJ�/�O�XHO��~�	���D��
C;>���ŧ�j
<a��NwSf~dP�j�x�n1(r��9*�=�mKy+�})#8����)���)�<(s�j�0$�_g>�x���)�$ g���M,_�#��q��/;��ɱ��T�5���ч�����9���������	�e飵?�]Y� ��o(�����M������<ߣ�ZW޸��m�3��[Lw||�Ռ6�}�Nw
�>GQ��5�3[���ck/����vF�܋�¿��v��� ��s5S~�z^\j���U
f����͢��t'����Z>%��Z�3�V�-+6bQ�)�Č�5��S���Z�iX�}]z�����u�Q�l�J��v��4(m�iՋ�hi����J:-�ȟm��F1�]?�0�en��K8��PuM����y\"�g�%lr�=n�q*�UѠ�?��~_�^\J#�l���&IL�x�W]�F0�
d�*�����p�>d�WgQ\e��)����"E��P˭� K_�	i����]��g���z�`�� Qp��J�D�A��Do羍���X΍��?~`�!�9��X��a��$ U
f����zyUC���t3���|M�V
))� q���:�&$�	I^���[�#D��mƥe/�0AF������<D4V�>�&�ȼ+��s���M,�#�;^p�{qB;��ڈn���p$�c��B���t&��w#>{�D�j���ɠE�xT{^r|:���ӥ
���C׹[%��2�`?-��W��|���]�xL��-)i�b�|��f^R����W���F��ּ�������J��pr�/�]��{��J*~?�OVt�[�w�0Q+z�r�K2��J�)ji�ڧJ <�,Fhh,�FY���q~��A�2�s�Z���<^p*:u�%S��'���G��R�߽���:�����\�M{�<�m%�[#К��v}�|��v�ݦ��5ny�Fw���,��AF�z����;UO�z��!�1���R�`YV_Q��d��pj@B�:��\�o\��^�&1�x�\t?�%vI
-5����7��I��at������� q�:��'*~r�6;P���le/K�����[�5'�N�G,������-���n���I�'l�=�����H�)W����{����.�(6��H�������-4	c�$bT�CP�԰��X�HG�~
T��~~������a�c�p׸%k� I�Rd�
�n�u��<�uF�i�`���FB��cj�U����*D�X�&���P�F��0��1�Y��<��e@$�����=�H�Q�n�q���o~L�ǡ��}����NO�]��
<A��$�@�]�JAN���(V|#�K�����;��;��J� �!���e�����\�g��-�1tS���ڰ%s��h\�4>�)��*����x�v�;�� v���}�qܙ���INv>z�w��R[h�7o�.)��ۤ陝�i��㷺��&I�Cd�����a��� "ZZ��̐*��@+�����^�6�g���;�tV���VP��n��p�?��n�������U�����_K������L
t!�!� ��l|}M��ۋ��� U��r��b��	��Ҧ��������t�jK��[�d��nQ���w
�V��V�,�2��R�~�j4��d:g��g(y4�5,-ŝ	*�F;��_[L
Cj��,��jql����¼r2�J�}����R�m1cw��ա�Kӌ�!�Z�e�|��kg��/ �"�� ���K��jT�=q!��U�qB��`��˛{�M)�t"��-��[4�40���q�7O���V�Gq+,�x�� �ž�'�a8Izd�4�[5�u9�գ�JR?��ﳉJ�y OܱT��N@��7Wܭ�T5��
�P��I(D�"��#�Ѯ�ӥi�)i���p*�O�ܓ	\#��h,���w_��|�qZ��
*�:"�Y��⎼pr�gp��K�1k���
b8����	O�& ����7!�FN��S�K�J�_����\R��|g�䪪X�{Z�g_�ywXS�%�a��{�@%%��Q�Ͽ�.~2Z�	s��2.Nl�{��
FL�ҵ�my�⁌e[6��SQ��C��i%zz�b��N-.~�ք1�wg�#;�Ǝ&�;�==�e#/��TVt�/�FF�����:r&#�U�9z�q�z  �������x�p�3�m����!F�ӶP���a}�.�`a0&<ш�$��I��~�)/�Z�����,���F\�H�bu!��ܼ���^}d��%��-�]*������5	`%س��:9�-y�߂Ⱦ�X��
B�����U�U��|;�ԁ�� �D$^"�~",�S�9 Z�"�$���#vpe�ɡwy�gc������|���Ƈc��C-j��ť7R��ٱOI�����CQ��%#�\�{�`�b��K��!7�F���,җ�+Mi��>������T�i�!�!t�Z䗂2�̕2�n*.X�A�/Ż4��l�&I��"E ��CZvgg8 �
�q
�u��'��Fh�@~�;񺞈b=��u vu�Gs$�5�H�
��5�LI��VŒj�\"Zn&�%�m̟0��&� �1�Y�v�������M����EQ��-e�#�)���n���xz��|O����Uϓ����c�!K�^�<�P��V]���V�#)��gh�ia,�	é���i�:}5�\�hgsC7�m���w'�͜�n��|��A3I/�k��<btP�8�m7x�/(��<�"�^�m�q�OR���>Y��=Z}o�<X��2W�l�s~�p3�������a,�yKJҢ���NzV��7��y��������W,\&��r�Q�&t�����S�]����kް�=�ww��W�2i�1�*
�;S;ݹ�Ѐ�S�l��-��6<tr&���oB �)�/����<�}�����Pެ��AH��/1O�ܩT�$9�#��8]��eC;%:�]r�)��ѝ�6�H����l�S|E~U��Y�Q
r[��į�^�mu<�����\�#C;�9�H��٣-�O�U�7������ �ԥ��1�_��EH̾^}�$2���-��vƚj/qNk���K8p�z��y.�;j������%&�f=�L��G$7yK�	��9w��H˄�W�K3O�ӞB(��F&������}��Gv�������I�:2���i3O�)��;�'�wy�8W+y�慺�x��B|S˃l�:E��E4ΓАÿ/vf�5���C�R�*y�k(X�r��4�����c�S�\)�)��sⅺ���J���qD��f�H�4��$�5u�Q�X�7���^V�38��[���[HrG��1$���K�c���H	���Z6a�ʗ.<��l��_U3� v���E ��2�;hM����
Xz�G�w�7��C����Du���@�M�$t��2��\3dk �7��_�-�5f�]���UC��`����7��{k�Px�TG��#�j���Vu�-1Ǒ�0�G�Z?LKX��́��)�S
dd|(O�zcM���f��^��ݬ�TP�	��]�r���p��e���.��
���pD�����)K�A��f��#��e؎^��C�e\���C�l�Z���γ��F2k9���x�C�?S��g�k�IFs�,�鐆c���.��@ ����$#n)`LQH�I!%hֺ2
TRXf�X�c�Сw:���]Ak��z�Ӎi�Z��8�$���XI�/�O�Z^m�����9���u9#�T,gJ�*w�f��i�u�Շ �d�ύ�|Wm����I��W��u��Q�LaMpF:\�4�hn<SY�����B�J���+�׹���!�-xb�W"��J�{H
!�^7Г�t\ژ�Cp�~Pp�����2nA��n,�a�O{���,��='���ܽU7y�n��l�d��}��+s�leT������zA�^�)�seU����eL:We��>�a�A��=���F��(؜\������#v�z�i�zy+ii|����`A��Sm�g�Z��XP��xg��2�Y��b9�����Ħ�}���󙯆�	 N��#]�Z�%�� ^�|7:K��O��XO��k�j����w��z����6����h����}K�Q����W����k�+L�.!�����P3� ���`\��.��1�����Ŋ�~��6��-�<��ـ�f	�����ow�2R����.�Nx�!��s"7Q#���(-���7șW�<�E��y\�}?�ޒ���^��N���0ٳ�_���\Si�d��3�n�7&�X	,��ɟ��P�);v~�=�b�y�89m�x��/8�F%�3����T�A&�){�
T�AzX�S�/Ѹ�=��#D�Q����I��'�f
̓m�v5��jD�j~�z�F�x���LtWg@�zz0Y�-��~���<t1cZ/����t��� ��:�K�C�^�I�; Za!���GI����O�Ƽ�Q_��h<�|�h��햇+b*7�l'�jQEq�+L4�l)nu|��B��`�U���j��{ߛ4�	,�?zd~E,@�N*��N(榵�pW�{{��rIM����땤���yT)������4ߢa��<rK#(�!?y[�Qg�F��{כ+��7y"-Oݣ"��A���e�pT��o3L|L?��Y/F⍉�7��BQ���t4qI�&k��lh۱�,�|?�^�S�QXdm��h�t�g��1�I�*�$0�6KƳ���Xs�߲���|ױ���𞊬 �%��"%��	���lg�4,W�?��k����-(H�cL��i5%��}��3R�{�pN9v��#�n�g�_�?'d�e�|�93�����>�>���r���E%��<�?Q��(��a4|1��ܟͲ��TZ0t���+�c/����@��)A#��Q�
�����+�� �`1N��X���C���<m4����!�!���u@�n��2�>Ӭ���9�גq^�D�)��_K��Ԣhy	6���9�	����׬�*����y}��f����!r��ԗ�VG��z٦��.�����j�����J��cZ��F�
HF�|�Vt�K��e'Ɯ�zb��:@%����|�V��pщ�K�E(�y�q΢�(�֮i�T�:�o���@��4k�yhTn|0���Cf����W<�;*��k$R�b�������׃(h�ܹ:)��2S�����1�=\[��ŀ�M�������6��Cc��_ʞg #yG���AK�@0�R�q ��t=�3}d�u�`��ș=6
���}�i�����4��!|X�A��9��!����>A���8 Ԉp����$(e&����"����`�M�#�T�x�D�C2���wٹ�' �=���]׈�`~����4�蔵���(N8���:��x�i�r{gB��>}v$��tR�ˈC����ZF���PG���-Ҥ&>��V���_^H�!jc�wkQ�_�@��%�$��2H)��;�6L�ᡟLNt���5��~7p���҄�H�nh�
ºH��E�;m��R�Î�Y�-����Y�+�?
���G�g.�,#�<h~��u�Bϱg���!��J���u�������j����~��ⲝZ��y��k�b���`���u�2)�Ў�)f��.�IF^ �q�'�݃R��m�E��RxC@����Gѱ�5�R%?¸t�� 2����We2l,�D�����~��^��o�qv&��<7�B璾���XB��N��������H����T��SBGF.R�3TSK(sNm$��>��==X����ag�~#/��B��J�0�D�/����/��!��B9�b�m,]�t�+���x�ۜ���-Z�W�g�y�$�^s�SB�y'ک[g�&5/�첍;$�0�9�屑~�\�*�[��0s���L�1M�׺�"g�_�4�"[�"{�C'���ON�aJ���IQԹ8��$u��!t��g�^.�#�@�S�����ƴK#����W0W\�$��w�1/�q�sK`	?D�>0��F���Jbd<���l���{��T{j��ʸ,b7�*݃���#Y��83w]Ur��4�w�(�z���{I�b���d��zǳ�!⻴	�tƲ��v�[��u�z��.}a�v'��{Oe�h;~�~ �Ƴ��f�&��X.!�آ+���@���r:ױi[ߎ��N�Jɘ����\�k���9�C ��͕}|��Ṗz�@��&X4>ƽ/�fU�3$f�P�=^YmU�hT�(-9��i-��ZΌ^����˙����	{7 ? e�Z�ܵ��$\���@3��R���q�x�`��@$���F��6��P�hJ�i���~@5�i���đ���-��
Y���f��4�*K��B�t������"7�uN&��j�[d���*�a�C08/�.�20f�d�#]`�o&,�;�|8�`�"�&Xi\u\��zV����~��1���S����g���+���t._B\o�UPH���v�ś��GxJ�fI�H�0�Y�ӷ]_^��������ީF'qI��;M�B
hÚ�S lR{�{\��H�,9ǡ��H�H��4�TY�0BI�yݝ�w��g�/,�d��s�(P��DP���d9�.���`�!_~��L�]ț����7R��'J\�_��,mwB�e?)uGzs��(��X���3p
h0��綎�FdsXh��˕�[�q�%M�
�$)h:��z�Jx@P�;��)^_<�{�L�.�CU�Ά��D:�����)LB���ђ/t��w������bR�d�T�}~�W���~r�/w�CY͜���V�(a�}'N���v�$#F�p�3����}Ÿ���sZ��R�g�k<�e?�u7ݚ��|@V��qN6q�r	Vy؏q�G��jqz�@��̊���iV�LYw�UW�~=��� TWR�LA��,g��C�� �����-=�H���_��_����)����X��7'��i%�;>|Tǹ�_�t"���v�	�o���j�[�d#���Z9V"1�E'A)���)
�mځt�gJ�@��'��@���k<QT�S&_ȫ��1��総��� �G��P������YfJB�yp�pײ���H;,`��U4�]��	��2��fBU$I5�N��Ȧ�N%N��k���	R~��e��E�L�k�<K8c�|o�6_,_{���ʿ�c�\z��'���=��ƨl`����GYy��=���Z��6q�\)�t{���=�4\���T��=��kq�I�w9,4Ml���K0ٌ��-�*��jOT�\�� �6�d���F�+Pk6��-�����d�e8�cs�ԫ ���\k��qʥ[�cf%��"����*�50T�j6k;Y8Ӓ�]��z���U�o3�������e��ICj��/D�1C,>&]��"�ޅ\�WL�X�*@�'�����W�b���H�aoX˃���܇t�M3h5ɽ��ԟ{�5).KFTY;(�9vx؄	T��8,����C$����h�D�'��|��<k$�jJ�N���P����4�\tz�b�l��e �@�ȳ�l�t�n���%VC!m5a{a�I�:�m��H7�еq_�Qb�2�o}K+�Ĥi�N�N}�}!˔��W����HR�V�����6+`���x/3�<�.g�K�}KZ:iM��>c���]�OF��������S��ا\����9���poIS:�n e^ ��)����`���k�0w= 7�ͭp��i��>�]��r��ކpü�����اf�m�v��0�����s���V�c��H^ ;� �l��1���i�Y���V>/c`hn���,�	�:����-kϵj "/e��Ɗ�Fr�N��pܯR纀0��V����p`T�d�4�Y!т��X�9���3:�N�T _
ա����tS�}UfV���� ����v���fKҽ�bxy��:��,����9����^�*�5��l�ߕm-$1�q�{ߴ�0�`$�($��T��)@�_�iIK�K6ҹ��~~V�J�Ԥ����^�ő�$/���?p��]߃<�o͌�=_���̋ͅ�:s���D��2��k�Z�
�T
/���|(H?�b��L-��2ղ�V#r.���'uo.��t'w���&����%��f;�\�R�� �Y�<�����~��?��_º�i�NxÀ�g\��W�FNmBH$2+Tѐ�N�4��D���  Wؘ̕��0l9����.�%�c�E�a��'��m�V�m�.��s��X�r�h+���f{���N�y��|<0���4����� ���N�!^3T'�����mN���P�>�2�ql}�c��z	���:g�
��dc�s͓�~���8�5�E;2�#���3}�#m)7�X�ʖ��m�Z����[������;%ۏ�̥��g*��}��-����7_�vp�ao[�E��+���ɮ���)<�F�Y�<>�t y����&q-��Rw��H��l|�<�xt����d��4։��O"@��ò�>𑥌Y����FLƞ�a���x��n���C��E:�1)��������s����5](��� tؑ:��\o�A��Y<�Q�G��$C�Y��G��vT�#{@����X��H��B��(��0�2�xXR��hĳC�_H�Q�dx�ʋS��S>���?�'4�B�`���(f6��߁��Fr�1���x�Ka��Cp�Re܍��˃��$X��2|u�8��O";[nOn7�oyΎ��I���{�8�k����>��+
�*���'S�K_�|��c?�h�BL�VL�wM'U�`vw�R||�^�?YRƸ_5O�����x���)Vȑ����h�˘S�����$���f�As0Z����qE�3�c9&�#�t��:1��nN����9�PAU(�Z��k�~���
�t;)���x2��C��)��p���=��+l�E�̞>ޠ��.��[2#��������:�T�Q�W�ţU��*�9͹�G��%�
z����/Y.��ܤs�K�����:�ѹN�w9�<ͯ�$�r���҆�ʛJ��G���SG`��_�M��>������-1e�\�f��V<��n,�>����[b�T��m-2���v�mx���:��u���=��/�j:��n+v�$���Q(�
� �����N�t��0�h���ͪ��1XV��wש.�<b�Dd�dL���v6t�b�?pEd<�.�QJ6�|�r�.H����C3{%�(R� &��r��-���(�}�a]��y>�v�ސ%�� �U�ۭ�F�S�����h��BNY�AjI��߳����1�O���\��U���A�hS=	���r;�3t��,|��3�r*a����Z�9�|J�Y����`$�1�I��]9nIpogl���|(�^�K'���F�妖��E�4���o������K^�xoS���Wkqx�싫��T�=((��ŘԣB�x� �[�o+5wo;����\�s�ҙ\��n��> Z� U��J��Ks˩�GR�C�ݛ��	��T��R�EawW�[,*�،ryoP�e/������-��Ʉ�ֆSN�Zm0{Y�%��Q�twQ`��qz�
�u�;�G���g�2l�O��=)��ɔTҐ�����9���FH@������$�s��o/�����\ϡob�Z)s�q�x�`_ ]l��,�coZ7H��G�=f�K?+���5���8Vj��ݐ��ӅJ�)�x:���z�݃Y���6s��9Vۋ3�^��L`�c��s_��t š�8��ޫ=�6�5�xA9�2�-�����\���8���� �ْy��=P��&���ы3�'�(m<��3HZo��s�llu��� HK�Q�,f���.}U��/��@��]�+*��
9H�Z&U�E�bӜ����H�I���u����o����8�����s_���q�E�z�	@�5���"����+jn �u�<+P���sm��Q��y�t$���$	�[����4^/��η�_&?��*9��rT�x�m�j�����Q��]r��Z)����`p���F��zЌː{V?X;3�R�==+}�(�v�U��=�¥	���ZF�~��S�_e1	D�1�8�°�[��p��
�A����T�*Q����+�V?p���T� =D�^����kܳ���`�b������(��ʯoen�N��S��M���c�#H�K4��8�.Lv֥E^���7��X}IJďC|����bX@��?�]΂�R�唢kB�����O����	����XR^ �S�Z;���'
��l&�nJp�}��]6/L�X��r��06S���=���7�#\/iH�S����Vg�Oc���
�X&[O=� >�R�M?�B�^���;0�KD(-�䊿>M����'��,_2�5����'��C�O3��G���È�-Ȑ���k�$��n��o�9O����>�fg�U=4Cɤ���e���hj`O� �%:[&��٣�0�>����t�o� ^N�Ң_#�ʜ�[w:=�\��� �0󟠾Ky]#x]ǁ�@�*�19u���@���Z��)�P������^��HD#Uw�!J�?_�`�9�c��ю!���̴;��[���/���ar���Pv������4�T
�Բe���Xo�p��JWY�ֲ����D��t+�b��b�vX:U���aI��O$�!���c���<l�}�@]�͵�#�|��#�N�|��j4��D�Qqh�?�������2i�snD�.���/����|�|#6��+o�Q��@Q���������q��R���=�	�8�l��l�p c�D1���g1
VP���$���D1K=�����|��h�0�����\��Z0S�DE7�'�Ea�n�&�G|I~2# [!&��_���_�Cfƪmy�8k�������άL }Q�Nq��˕�����g*�R�p
�U�,�n��:>��hx�}�)��&��|
�g�y�q��L��qt�mn,{����\��j�$I/�P������x��Zh9�ج�K� �T?~oQ3g��1t&H��{���/_��\�B�H����_��~��=����?cJq7�D@Q�b�B��}(�SL�6T8���|��� 	��#��rkڦ���L(M��4�����a�O'2(������S��)�a�����8p�������	+8��oF��YLw�2��-8q�v��`22���)�XK ��X|i�w&IZ�=��][�[�ށ��*�L��h�7$������=���N�8�ݨ�L^�7 4�.lq�"�#B5^EϤ�?��i�r�J�[*\w��l?�MXi��SG�@gZ΄IFA3VfZ,�����ٺ~B4�e2�5��V��z�~�́��d�D�c]�o�?u��(���Zd����96=��F/6���>%��Z��p�-�@O�1��E��Y-�go�)S�n�J<E&h���̉)'v5��[� �~�j��G(*�*�s��3a7qR?-G�4,��۽�VnV곰j��Y>i�&n���pc[�׌i4��=�(2p��+�V�Y��։��_Fa,H�W��w(k��8���� �D��`��0c���$NK%9|��7]$E�J3�:�<}�?OE9R� D��:	F�S)��*����;����I8��C��87�3z�m�&�pO�{�����.���OEV�
w&�p�ԉ��-��꣡f�
6�
�#J��+��pPh�
���F�O���,��U*n���Y]V���fD��A�JF�*��iV�l �m����50�\��(jxu�`!�p�,��9y� 2����ֈ�'������r ���|
4$GM�j���KJ�fFp1��̓āׇ<����ëd[��s0�Zh|ڸ"#�� t����K�x�|�Z���m�m�xJ|�`��=���kq}��׼XE�t�~�lW���R���
.��5�B�����&4���u��O��m�a1��B�̙��-&�l�Ԩ�p���4zIw&�v<Pz�[Q���A-��ݸ�Yж��gP��;��RJcSl*͢��E:�t$4�]/�x�r�S�RP�����L$֑�����]���CjB�=�=[�PQʰ�S��X���K�ۏ'թ��g9*�k�!�0�Kamui�!�e\��iz�����8C17�f ��0�y�����|�8B��?I��32���U[3�A�}�L�?�M�2�������΂�U�T�x,p:�w�ԣ)�܅��{��ւ�S��A��$3j�Q�~��!AN,��C�B1�mV*{�蝝�i�v�"��H%S���7��߃d�*��-���;~E3��󞣧�M�7�����c�*DT�3��謽.߭q�U��8'���^�}0��|Yi��hԉR!M8S+-����EW)	=����,�B�ǀ� ^X��xS�J�Y��^>�^�u�O�|�R���b0�EИWX+�n�x=f1���d��G3ʓj��6\2�y�{�3�؇H��"=�g��Ո��{[)�Μ��x
�08��v(�)�6�>�-�����w���Z�z�&�����t<h745�.ϛl܅��vİC�r���v�pȦ��_i��oLY���hq�yȯYkh�g~@�Lv�ö��þ�Ɲ���M��u���<��`�]�nu�ȭU�)��(�R��8�������>,�'zDʉu��Sv��7�S���s�����d�/����}f�/�Z�#��Ø��U�J�]�LokB�=C���ؤ�6uk�;Eq(e
�����#�N��tn��BU�;-r&��a�P�ۧ��IfG1�؂���NRYꡓ`2G�1���3��>�ҫ�T�^���;
o0b[�Z����M[��Gl��5��N��P䢫z��)�f3]Nc���^�iS�ѝ�����#<�'F��k����;��#'\s�ZA��%����w����t�z{���c��,�謯���) W+G�?Bo��.��$`�@!�5���!|n�Z�e��#@�*�rS�U��/�5�e���$��p�%�%��r�F9��2݊J|tֲg$�k��O�[�p�Wo�;IE!�#�T��9��D"|��S����G�����כO{q;VZG�����A ��tZ���J> ��~������̋�N*���������1���J�Z�q�P�'��l��Gƫ����S�yq��|�z'ta�Vw�Id)�0M��|��ǹm�<���l`CD�5
�q�8J���|`�c����r`{�-m���t餺���:����PD_��8���/��aF�Uƣw��倂�tMs�*���r�V�"ƺT\�fb틀��E�F�O5u�Or�1 ��\�����v9��
Ǖq_�@ �C�Ra��ʆ�����2�k�9��]67yO\�+R0��&��voN�#D/����OC��.N�t_��F|*&��~J= X|���?G�;y�)�
J�b�I�� �dѢ���� !��X��l
B3����DD{=F��d�o��AF=_f�vq�F����CdoVl�Y��$Jb ?3~6C_�]���'�7G�Vg9c��k�)��r���8���o��pDn��$�k$�	$O7�L��Z'F�/ �ȽXo�9����B�@*����>��\�C|	[�$���/Ft5�Ԇ�����^�:���o��U*&w1O:�҂xy��/��=��v�mp�:J�#�F �gvD�l��ܡ���<�Wp���n �'�l��b1���bR��X$48�*�埫mE�l����:$TF����c��Cu�Q>[I�F�z��m�;;16VfCp� ��ܨ��Q"�����U�[E0�AG��֙-��be�(%'���Fk H�o@���`��i�jlĶ*
c��6d~�������P﨟S��svEcg�%xcPյg�$��oжiC:b�9�3X�nɛSa���qZ%����p6�֝�+1&�Jd�|:���\^V1{�kh�c���h��Z	���2J[���ҖD��]�K��G!������ӥ&�n��ؘ�RPx�%�U�Re��C׶�Ӡ�l���<Y��Ɂ ��"����gI�|��e��IP�Ѫ�{4όb�H~9�ui<��$F2�|A$�߯��í�ë{���SZUt��/�ܭ�,��64ѧ1JY�8{��;n[|�N}�H/��&�C��\u�<�$���ׂ �bFt-\˷�yE/"�*�8���x;o�7�Zt𻐻��h�� ��>�d�'���7x[(�p3��u��꘻��֞{=�.��ѵ��H}ᐏ��>�.���gqU��f�k���@��k��ô��A��W��z�9'P{t4�@�.�j���ff��0����[�q-P��M�Dp�u�#��s"�w/�+�Q黣o͔(P40y�AP4�%�
�����ڊVfg�j��Af�{������p��֜腊���q7��K*���K�),�#k�7	�@�\2w��஽�2ȢM{�Sa�"![C�ŷ�Tl�F)臩A���M��j��9\H��p�0�݊�}4��O
��!HZw���o���e��:5d-����7	��T��J�2�՛ZDL�� )�����������P��D�Hn�:��bK��^��!I����		���B����J��|pz���|��4����$,VUB����) E[�(Z��V9�	E1���	���IQ�&�c:�1�Z�-��pj9�Ty��#$��2���	��kԯ| dRj%34��Zګs#pK�?�y��UG�6�i�`.[�4���5��L.���tnI%߄/Y�y����N[*���Ah,����6��Gq<������%.Ւ �(;�2}�V���_2L��7*�ʌ����@�T�;����;�y<n�Հ(�ƀPɣhX�͉Ϫ�k�&�ճ�wQ���⦶�I5#�6��n��s�FLޙ�S1�$�fc���R��c��O����|ܯ� ��]iI��m�*��5g�K|��;t9�S$Z�����֤2���su��ӄ��W<�d�1�F~��1=�'7*�4@>�u
?��7���8L��K�/-��[>�����e�_CI�\,Iz[��f�j31t��� ��q0�	�u�SrE����1��$�.Jh���y&.���F�T3@��*Dņ�l�E�IJ3_� ?J3Իk�|���a�w��^�����N�bp!�r��i���s+��T�G���P�F�/RQ�r�o�_�m[��
E'UlRt� �z��u��"�O��8��5W|#D�Jz�" ����z5��|;�Χ��>�mk�����S���K���[Y�̔8u���7!]-��R�L9 ��4d�����:�'ZƸR)�Bd%�c/& F��zp7�H����՘���3\B��mᣃ�.�ACF�R�AI?Bȉ���s�����-w7V�$��wǹ���Sc��L�=��A������ڝ�E!6ɡ��ˏ�sS� ��m陵���p��n�)�㰉U�n0�IWp����˓�����^��0 v#��{j�M�[fл7h���+8�(XVb��_�נ5g�0,Z���
��_���x�NSNtL����Lw��JM�>��۾Θ �J6�,S��e�%*��pW;����Pػ�(�c�襲�lc������U�>9Eg S1Ṟ=틢���=���N��/��z��������F�2�	�l�G����3/ x���_�D�p�na���Q������J�:�]P��ܲ L�(i!��J�G��e%������J;��-)��$ۡm��۾.�t[qR�16Y*�du6L)���9�p�t���n��!;��B���y�]���Z00:A9z�.*��v�ZI����U=b����<ϸ�崃���.=e�[�.�vi��[��Jz~���*8���@��]�]��u7Q����f 1�S�wb��'a�=�e*H�Ϥ�M�}�7�������y��P&�5����ǫ��U���w�j^Vo���% �{6�6�h��h���9�r�v��?1��fN������ 
-�CO<X�I��.�ԺA�$k�1x�o�p�VٟB�}%GW�њ�V5.��9\�{&x����$C"g��zK�a��:l�s�:���2��F����F�էcQ]�RS-��V`�A1������А�4�?�$�>4gy�y�Hn��],z��ܽ�2葦,���y�8q�|�U�i����J@/Z�N"DT�YB�{>�ϫS�ˇ�U�4�@O3����6�S��!���a���l��x�<>�����,�釳v�_�hˇǖ�N����o�ljmM�R|b�����T�������߼�:I�<ZK�KÂ�����4��c�|�������ON)�w���b����:R���[P����a\+��5٥�ߜM��K`H�=}�rG���'�r�NW�u���R�C1N�)��>y���98�tZ>�H���>�T�5F3D��%���4��Qϼ�%��C��>N����+����a�G�������m3�T�~�������`yy%"JS=#D����{oXU�P�P+�x�a�8�;����������+�]��ϱ�p�-���i1ϼ����\�����#粱0���.l�5r�y~$�8��9 sڟ��V�xh�f�W��
eMY&?�s�m�tl�]�H8.ɹH�h���#�y̸���%��CH8�Jx؋(pב��gpq�QBn$D�`�� ���:b�A�o����MT���A�MML��ڲ�'��k�FfҞm@/\Q�$��B0���b����,��s�7fR"�0o�3xY�S0�Z��6�t���:��5����<�L@���p0�b�8�4M1�wCG]����~\��񈻲��&?-@!�� ��gA$=F*9s�� ����P�QO��B��?-2t$�f���#�
�80h)�`�-<��A�	�wO,@w����J�]}X1?j������c��R�L�&���kG��Uc9P������j.[֡����)���٫~���$`��5<Ds�В^�E�da�C�s��:]�Q�
4�D�f������<��|����\:�}���E��K����
�Ӑk��)g��x�����W������c��2B]/S5P��t�i�����a�� kZB�0>�Jw�=��~��Cf�U�vp�+d`uzG��F���*�vI���L���:�c'����%����?
��ǫ�&�d+p��,;���h��(m����8%:��)4
�d}��RO���j�f��g96ؼ�z�	��<m3X��R�uۜL8��Ip�c���r�L`vl/��X50'�v��^E����j�>}���?	�1X�� �[!������ȴ�|�[T��8KZ�f�>d���qt��[�l�=��/���1���d:X�����_�Ϊ=�R_�B��2����h�S�!|�����F�g!�Sq�+a �- ft���<��V`Ƙ�"�f1j1&�n�ѫ%���p�c��ut�/1�b��J|��J߰�S������������T#���/�!��E2��7S�*'r~�R���Ǚ�*!$�r.����_�ts��u�`ݪ�����1�S�&���gꂼs{a�.��ǫ�_$O{���� �\�T��tsЕ���,n,�m��pOұ���XF��yP�稸��-Ng܄Q�]W4�j >��\��縔���JU�~�qsY��8�#�vt�Jve��ֱ���HW6�I���x���v�����CI�w惄�W��b��AsLMDQ�>��DѲjf���2OU���%(�-�i����t��jeK��W�,��$&o6$F���is΃��J�}��#��B���E��
8��[������ѫ�L6*
H���ɹ����]F�FN�?��5H����m��Zc��*"�r�I,�P������ܐH\l�'#ܯڸ;b�C5�v�����j�����$j�U�x]��O�^+�����R�>R��h\��Θ��l-��l�P$$r])�ţ��	S,�7�N>� _�|�f�*��JoȦL6��|ܻ�#�!D]LQE�]�-~��
~yŒ_)�� �����{�*n�������M,|A� b���;�,�DB&s���)�i΅nh/��� f��`<Z�������3^�O݃���dyEQrB�r��O�����k�H��5?��m�{�# 9�w��j�~
-�c�1�ƈ'6��PO�5׾�+|����� � P?,6ob�k�(�;�&Jڒ|Z�`Nh���ߡ��[{���b�ʩ-A2��G�ZX���f��{?��6����ͯ+�Q]�s�����h���b��R��>�{���R�UĘ(�tg+�Ą��Œ7�����ߦ�$&�/	�[GP���
�[�N�������u�"9kt���|I5aVĽ@�c
]�j�\(b��xfz�?���+�2Z�q����r�`��+�:�2z3աT �M�bC�[���lX�wڧ��b���(\��{�n��־oϺ2XC�Ra�Î��p:��,3�U�IP�9#$�x��M�1fg�	
�<�%�d�'��.(���Mp}��J�eK��5aW��M�L6�؃��X�(��|���=_c}a'"9x��`֊�k�����@�+K�ΘT���z��@����(.�j~����XofiN��Cr&�Mn�&,Y�6A��8T����O�T�"�#�7"���h�	��m���y{ޱ���v&4�m�!���MN6d.$�"���j�f�8z�쬄�)�s\��}��}�Y�B�2Q
���= ����t��>�3�q�ig���%H�#�,q����� 7�}]��J��CN��?Kj1�vy�[
nV�4}�VN`�\0ʞ�P�CDN�jQоR��bn:]ϝ� �t���0�|	�	N CC�b��Y�+�����ihGSKOjµS#�L��^P#�`.���y�ΝEu��'/�6�ew��U���!V
��44Μ�,ަ�T��{tDw�g�6X��\�0 �k���3lA짫�מ֝��J�O�q\�M |��m�{n���(#�^�����܃��F?EA����0|8lW��Ӱ��$au����k�vk�$h�Z��W���cv��`�֌^Z�=ڶQ~\���ǌ�h�
PK�r�������?�����̾�d�S��L�(M��Ń%+�zEEM��7�ۧ+�*����f�D)fT�q��u�9������q|i��\ j~��.���'���{K	S�ނ��+�}�G��h<�J֝�������w���@��t!��ẅ��&��l�%�Hl�c�����L��j�D�G;<9K+*�V��
�,X� vv�Q�r<�����ہ}�	J��+lx����i*	�PS$�560Z���}��1a��.n�����3o�6���%Nm�&m�.�k2���pb]G���� 8=Z������t���M�~[�����h:�X �~��rC�-��3A9,�>���U����ȝ�k=Q�-[�d1|YY
}��0�?����vM��a�Q��Ms c�XA�M�dQL2l�5��D+��\�/�{k9M�m�|CY���M�,o1B�j�΁]ﲟ�Q��2�}NK�f�"���|rޜ�T-$y,�a �W�i�Z��~����m��Y��Qp�w������Zy�D)��.� K�;�^�έZ��D:j�I�/+d��J]��R��%2ñq�����1�>ᩈ�{���\9����:�[V�s�$n��c�2
>��=�4RsZ� �uP�B�?����yR�V?[��������VeH+�TEt��h���7�2y��)��PJ�Tϩ�A��j/�N�載���^&ȳ�<��¸�]�w!������][Ʌ ��7O�a 
f[��"~�(X'�;����f�ai�Gk
�f�٠�(�i�X��	�!3��K��Z>ᄴ5-�ן�~��p�@�d�g���ő���A�ΙQ�XUx7Hrl�U�z�3�	���
 !�F�ڲ	�phbU��^}�<�{�\f��W�{Im�8�JQ��B`��"���α�"m"����x����}Э_W���R)�ԩ0WG\7�g�u �s��Y��DS���^n�#%>��������T�Us���&\Bt�
?�>�єC<D�&J}�u����<��q}���PHx2����(2{���Wt�׈a��Iح�F�L1�X^X�C``���6���>���ܸ���5x��z�"ݼ5k��e3"�
-��zs<����d�`�/qC�P�u���"�/���$�I�����~�rڛ �$(��g{�����
��͵�?]@ܦs�Ic#+f"�}O���.3u�0k$��qq�׋�Ң��x<�>����y�HZ���ſ@;�Xp���Lhb&�Sql#��Q�Z*z%�d~p�O�ֻ~5����=ǧ�)���$������!��^ƒ%>觢F��u�	q����c����r����D��a���^&o2p�R��2������%´�;��w��'��۪��bs��Ok���[��!������
2p�܄���ɨ�'��Y�|��:T޻,���:��EmG���A���	��9�.{x��c�\S�f>\���u��a~���2��gh�wT��� x�/+��O�i�M���#sW#|�N���t&ᤣ�����,Z࣒��NҌhv���k<r�wI��u  Z����%�wV�����faz�R��H�)��2��UU܍��&Z�[´��PH��c�,W����Ω$������8�w�BM����`W@c"�����Qj��ku?S��`S�«r5 `w/�Үa9]x"إ��%a��,��Z����Sp�g#1pa������ҹ{��9���py�b&.�6��d@E �h՘�{"4�~�sx�s	���[p� u���4xF�Vt/�����n-q���h�`
��"���pHf�W:����!,�Z
�E����[�?�$K���O(�����~/��0��/a����$�k3s�4@��[��@]4���A^P}%C�uı�qf�͛^�6�B4����hW���I�Z�f�� v�H�3��6�9u��Vi�6'&�x�����ۼi��~К��X6����T����N�~�3�S���)������.�ʶ�q��[ɆeJ(��<�1�nd�9ݔR8�F��Y�{�,Y�6�}�ZI@��rL����$e�O1��_�luX���c�h����솉�5LD�3�l�.$�(�k�]'b
�İ�TQ�Q�J6ohbq�H�P#b��I��}����ǁ�p�:NE�oe��D紲w�(��n�"�M���QB��|zT$����"�6މq�F5L��;h�]����Sd�g+��v���#�y~l��۽��C��Ҕ��G�g�G�'|��/�y������ͮPoF�_ULI��W�tE�pB��*��;)�Rse;y'm\.`�P��p�A�y����$��j�Z����#Ò���&�����_���ޣ̃R e+僩}��m/Kᕮ��{g�6�XL�Q���}�&"���Y�Ҟ��_��k���{���vr���o����aN*Z7��C/��J�O�@����������B	�Α0)�V�� ��&N���L�T'���|9�&�N`�#*S�[�e���-*�N���p!N�K_(ai�WcNc��}RH��C~���L�I�ɿ��>sį��װ9*�"6d� �+�hĞQ�l��`��PTp��Cb�fS��g�u~��Һd��a�<��[����d�����D�g���� !��?^t1�yԚW�zRݽ�x-T��\q�ҭHk�e�9�Y�{jvM��ȎP�o�K\��lc/�����^�Pzam֓�ބ�4���!�^Գ?4�,Y�ҙ�y��]�^�Ǣ@bA��0aX�F|k�P�c�u�&���S0�@]��ܛI��t��J0�vm^F�&�'c���J?����+g/���t��+_i�g�a��z}��w�U�;9}=[E ��?����W��B�bx�eЏ�W���"՝�T�tG�b�a�Q �A��RνqW22�2ҁ][l�����a�S���h���&Y�t�yZ�ΊրB��+�<@�`�~H��q�q� 35�q��L��8�ӝ�{�w5���b�Mj��-j�ePrz�e����^EE����٬?�<�q�B�ʻ���*^�O���~�{#p�)W�^K�:��}��vǌ���v��٦�n�/.S3�ž2�A9:���$�X��"�Һ���w.�jy�"����0�X�I+If�F�O�����7��b���p�g�g����n�g�D萄�mGԝېETe�,�hj˛����GZ�c��ƫ+�碭w��4y~dv�N�0fi?�K�(��Fj֮�v��IR*�(*�?~�X,�s^���ϸ�f�'����V=�����l>s�acR��+�/#c�N�\���%�[c�QQ�Ktꆆ���� ��Ov8��-.�I�I��N���G(EÙ�u�sU�vB)�'�s)U����t|���	eN90G� ���&m|Z�M%@��LW\gG��8����"l)��f(�**R>rW��~S4s຋6*t�+שلh��=������Oe�2�v�����"��D�~�o��*��m<JY�-2�5�W�s'L�t?��!²�$��'���ņ�Mf*C۷g��!�����r��	����Z��~ɭ��u�@�w��L8Ӈr�#��4�v"�HG���8��˲H�  �Iښ�&�4�h�&_"�D���S������ 8I��x0�q�3��.������g�<�~ku�cߥ��<}�O˺�ܜx���O�2���D�Q-��ֺ˂c�-�*����ė�W]X�A��	��1v����N��P�яa���e��aT��b~�r8��S�>�}4B��n%"���
d�\*�nP�f�g҇��
Q#��\����hoP���Y)F:�,������8O�/�TE�� <N�~Q���^���/�G�$���7馏�k'�rk�(�׽�O��r
d,�.�`#Bp�oJ��3t��������W5jm�u���JW��'ON�Y�׵���O]��!�"5�Z��?���ȷ�R�{�
޳�����e��\	��=l�2F�
�S�k�F�	�T�J�u���3Wg-�|�\��]����2�D����3�k�'����xfZ�:�|C�om���v��h��%d������{W��?#u��gJ{#��բtY1�6��U�ᇧu���LAo_/"ݴ�pT�":w�K�.�v�}9���Qþǖ��DwQhǛ����`O�_4&R�+`����Ls(��׬�|6 ӹ��.'�EqL���7��zq���&�������Kht�b���c����p7���*��yk��0Ɩ��!,Bm����-�|��F���f6�����O�U��d��lZ�ϣ���ode�4>.;oe+Nq߅)��WK����Y�����*AB���F�|�L��$��n�_h�m��F�F����9PǍ2>c��Q֠ *C�ߠO��1���O*�X@��:�;4L��P�	{˒�K҃��Q����b�7�4rR�*��A���1}�a˯�%�v�� ��0B�@?�<���;��L��
7K�*���T9v}g;
kd)1r�Y�8V��JO�����Ԑ�h��(S�O��M��k:<Տ��_ܠʶ�ٳZc�J�|��T�M����|�O�|��k斧�򥇌�@;�c�X)2 ��ʬ�G��M�-���F6h���d���5�_���k���T1k����718�@ .�R�4��[��-��^��[ta�%�"$��oZH��K�6W���$�9�H��6e-\�K/��a@.��X�j������m��O�F�����Hu�o����@�$���\�I�{�^\j��b��%]l��Ռ��j���r��=���3���ɿ(���K_�$�����oM�#�X��(Bi���I�_q���lJ'����w[�.�%f$#�Dg��7��8cA�f�$�O)��G�6*i���К>��X�cJ��
cZ��	��~�iqmZ�(Ȯ+�J���G�5�6�o=�����U"�O�u�?�����f�־J��N�;�lR�f�z
\,��+W�I�4�<M��<��k�o<���D;w2K,T�0"�\3��'Cv5#o�mA���J�����T�8d��w�߉,�}��D�:_zὑ(u�Ց�xT���%�����i�È�f��R}���p�o7�B1Zh�x,$?
q�����Ʒ�xσ�\ �&�h�Ԉ"Bj��)� ��!8L6ǖ>Q�GV*Y�,.��[�ϯ�j�j��OZ�=]B�:L�B�ً����s.��=e�#�v\���NZT�?��>[���M'�BJxn�+83`��I����o`N�'�ZG�'���U�ՄX]�W�oG�����7᳃u\Q�ޥ��WXg�w|<Z�4�Rd�U�+� �M���k4C�Ұ� uw�6}+��mce��k#��Zɰ.9���Nɓ6��3��,�^�" �'J�.!h�<��BJ�@;x� <�0�.T����.K�Gvy�������9�O��L�#��˔�)S)q@Ӎ-ц��,�L ��[�O��ڃ���5�֘��w��~�_/)v6����B�y��҈c5r��_wc?��4���3�]�w�PS4=�fY0���/������G>��w�ia��ew䪝t���ڼ�bL9%Cg��Xa	]J#��OIs҉�M0�l�F7HLX1�"#�~g��&�8ݽsOT-��-I"ɡ�2Ӊ j��{�ު��w�|���{����"W��m!��C!���t੬Ɖdu�Lk/{f��{Y�v��m��/W������IS���P%%';�w\DW�la��^���ل�Tٗn.���ڵ�[��рG���$����K,��6��˙����n��n""�j��-�������